----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 			sergio rivera (srivera (at) ucm.es)
-- 
-- Create Date:    	16:08:08 03/02/2017 
-- Design Name: 
-- Module Name:    	histogram1024 - testbench 
-- Project Name: 
-- Target Devices: 
-- Tool versions:  	
-- Description: 		this HW accepts a binary pulse as input
--							and classifieds it by its time duration
--							in a 1024 bins histogram
--
--							it uses 64bit counters
--
--							the output cable "hist"
--							is the serialized histogram
--
--							the time resolution is T(clk)/2
--							as well as the time base
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments:   this is an initial version
--
----------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
  
ENTITY histogram1024_tb IS
END histogram1024_tb;
 
ARCHITECTURE behavior OF histogram1024_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT histogram
    PORT(
         clk : IN  std_logic;
         rst : IN  std_logic;
         Pin : IN  std_logic;
         delta : IN  std_logic_vector(63 downto 0);
         Pout : OUT  std_logic;
         total_time : OUT  std_logic_vector(63 downto 0);
         hist : OUT  std_logic_vector(32767 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal rst : std_logic := '0';
   signal Pin : std_logic := '0';
   signal delta : std_logic_vector(63 downto 0) := (others => '0');

 	--Outputs
   signal Pout : std_logic;
   signal total_time : std_logic_vector(63 downto 0);
   signal hist : std_logic_vector(32767 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: histogram PORT MAP (
          clk => clk,
          rst => rst,
          Pin => Pin,
          delta => delta,
          Pout => Pout,
          total_time => total_time,
          hist => hist
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 
   Pin_process :process
   begin
Pin <= '0'; wait for clk_period*1/2; Pin <= '1'; wait for clk_period*1/2;
Pin <= '0'; wait for clk_period*3/2; Pin <= '1'; wait for clk_period*3/2;
Pin <= '0'; wait for clk_period*4/2; Pin <= '1'; wait for clk_period*4/2;
Pin <= '0'; wait for clk_period*5/2; Pin <= '1'; wait for clk_period*5/2;
Pin <= '0'; wait for clk_period*6/2; Pin <= '1'; wait for clk_period*6/2;
Pin <= '0'; wait for clk_period*7/2; Pin <= '1'; wait for clk_period*7/2;
Pin <= '0'; wait for clk_period*8/2; Pin <= '1'; wait for clk_period*8/2;
Pin <= '0'; wait for clk_period*9/2; Pin <= '1'; wait for clk_period*9/2;
Pin <= '0'; wait for clk_period*10/2; Pin <= '1'; wait for clk_period*10/2;
Pin <= '0'; wait for clk_period*11/2; Pin <= '1'; wait for clk_period*11/2;
Pin <= '0'; wait for clk_period*12/2; Pin <= '1'; wait for clk_period*12/2;
Pin <= '0'; wait for clk_period*13/2; Pin <= '1'; wait for clk_period*13/2;
Pin <= '0'; wait for clk_period*14/2; Pin <= '1'; wait for clk_period*14/2;
Pin <= '0'; wait for clk_period*15/2; Pin <= '1'; wait for clk_period*15/2;
Pin <= '0'; wait for clk_period*16/2; Pin <= '1'; wait for clk_period*16/2;
Pin <= '0'; wait for clk_period*17/2; Pin <= '1'; wait for clk_period*17/2;
Pin <= '0'; wait for clk_period*18/2; Pin <= '1'; wait for clk_period*18/2;
Pin <= '0'; wait for clk_period*19/2; Pin <= '1'; wait for clk_period*19/2;
Pin <= '0'; wait for clk_period*20/2; Pin <= '1'; wait for clk_period*20/2;
Pin <= '0'; wait for clk_period*21/2; Pin <= '1'; wait for clk_period*21/2;
Pin <= '0'; wait for clk_period*22/2; Pin <= '1'; wait for clk_period*22/2;
Pin <= '0'; wait for clk_period*23/2; Pin <= '1'; wait for clk_period*23/2;
Pin <= '0'; wait for clk_period*24/2; Pin <= '1'; wait for clk_period*24/2;
Pin <= '0'; wait for clk_period*25/2; Pin <= '1'; wait for clk_period*25/2;
Pin <= '0'; wait for clk_period*26/2; Pin <= '1'; wait for clk_period*26/2;
Pin <= '0'; wait for clk_period*27/2; Pin <= '1'; wait for clk_period*27/2;
Pin <= '0'; wait for clk_period*28/2; Pin <= '1'; wait for clk_period*28/2;
Pin <= '0'; wait for clk_period*29/2; Pin <= '1'; wait for clk_period*29/2;
Pin <= '0'; wait for clk_period*30/2; Pin <= '1'; wait for clk_period*30/2;
Pin <= '0'; wait for clk_period*31/2; Pin <= '1'; wait for clk_period*31/2;
Pin <= '0'; wait for clk_period*32/2; Pin <= '1'; wait for clk_period*32/2;
Pin <= '0'; wait for clk_period*33/2; Pin <= '1'; wait for clk_period*33/2;
Pin <= '0'; wait for clk_period*34/2; Pin <= '1'; wait for clk_period*34/2;
Pin <= '0'; wait for clk_period*35/2; Pin <= '1'; wait for clk_period*35/2;
Pin <= '0'; wait for clk_period*36/2; Pin <= '1'; wait for clk_period*36/2;
Pin <= '0'; wait for clk_period*37/2; Pin <= '1'; wait for clk_period*37/2;
Pin <= '0'; wait for clk_period*38/2; Pin <= '1'; wait for clk_period*38/2;
Pin <= '0'; wait for clk_period*39/2; Pin <= '1'; wait for clk_period*39/2;
Pin <= '0'; wait for clk_period*40/2; Pin <= '1'; wait for clk_period*40/2;
Pin <= '0'; wait for clk_period*41/2; Pin <= '1'; wait for clk_period*41/2;
Pin <= '0'; wait for clk_period*42/2; Pin <= '1'; wait for clk_period*42/2;
Pin <= '0'; wait for clk_period*43/2; Pin <= '1'; wait for clk_period*43/2;
Pin <= '0'; wait for clk_period*44/2; Pin <= '1'; wait for clk_period*44/2;
Pin <= '0'; wait for clk_period*45/2; Pin <= '1'; wait for clk_period*45/2;
Pin <= '0'; wait for clk_period*46/2; Pin <= '1'; wait for clk_period*46/2;
Pin <= '0'; wait for clk_period*47/2; Pin <= '1'; wait for clk_period*47/2;
Pin <= '0'; wait for clk_period*48/2; Pin <= '1'; wait for clk_period*48/2;
Pin <= '0'; wait for clk_period*49/2; Pin <= '1'; wait for clk_period*49/2;
Pin <= '0'; wait for clk_period*50/2; Pin <= '1'; wait for clk_period*50/2;
Pin <= '0'; wait for clk_period*51/2; Pin <= '1'; wait for clk_period*51/2;
Pin <= '0'; wait for clk_period*52/2; Pin <= '1'; wait for clk_period*52/2;
Pin <= '0'; wait for clk_period*53/2; Pin <= '1'; wait for clk_period*53/2;
Pin <= '0'; wait for clk_period*54/2; Pin <= '1'; wait for clk_period*54/2;
Pin <= '0'; wait for clk_period*55/2; Pin <= '1'; wait for clk_period*55/2;
Pin <= '0'; wait for clk_period*56/2; Pin <= '1'; wait for clk_period*56/2;
Pin <= '0'; wait for clk_period*57/2; Pin <= '1'; wait for clk_period*57/2;
Pin <= '0'; wait for clk_period*58/2; Pin <= '1'; wait for clk_period*58/2;
Pin <= '0'; wait for clk_period*59/2; Pin <= '1'; wait for clk_period*59/2;
Pin <= '0'; wait for clk_period*60/2; Pin <= '1'; wait for clk_period*60/2;
Pin <= '0'; wait for clk_period*61/2; Pin <= '1'; wait for clk_period*61/2;
Pin <= '0'; wait for clk_period*62/2; Pin <= '1'; wait for clk_period*62/2;
Pin <= '0'; wait for clk_period*63/2; Pin <= '1'; wait for clk_period*63/2;
Pin <= '0'; wait for clk_period*64/2; Pin <= '1'; wait for clk_period*64/2;
Pin <= '0'; wait for clk_period*65/2; Pin <= '1'; wait for clk_period*65/2;
Pin <= '0'; wait for clk_period*66/2; Pin <= '1'; wait for clk_period*66/2;
Pin <= '0'; wait for clk_period*67/2; Pin <= '1'; wait for clk_period*67/2;
Pin <= '0'; wait for clk_period*68/2; Pin <= '1'; wait for clk_period*68/2;
Pin <= '0'; wait for clk_period*69/2; Pin <= '1'; wait for clk_period*69/2;
Pin <= '0'; wait for clk_period*70/2; Pin <= '1'; wait for clk_period*70/2;
Pin <= '0'; wait for clk_period*71/2; Pin <= '1'; wait for clk_period*71/2;
Pin <= '0'; wait for clk_period*72/2; Pin <= '1'; wait for clk_period*72/2;
Pin <= '0'; wait for clk_period*73/2; Pin <= '1'; wait for clk_period*73/2;
Pin <= '0'; wait for clk_period*74/2; Pin <= '1'; wait for clk_period*74/2;
Pin <= '0'; wait for clk_period*75/2; Pin <= '1'; wait for clk_period*75/2;
Pin <= '0'; wait for clk_period*76/2; Pin <= '1'; wait for clk_period*76/2;
Pin <= '0'; wait for clk_period*77/2; Pin <= '1'; wait for clk_period*77/2;
Pin <= '0'; wait for clk_period*78/2; Pin <= '1'; wait for clk_period*78/2;
Pin <= '0'; wait for clk_period*79/2; Pin <= '1'; wait for clk_period*79/2;
Pin <= '0'; wait for clk_period*80/2; Pin <= '1'; wait for clk_period*80/2;
Pin <= '0'; wait for clk_period*81/2; Pin <= '1'; wait for clk_period*81/2;
Pin <= '0'; wait for clk_period*82/2; Pin <= '1'; wait for clk_period*82/2;
Pin <= '0'; wait for clk_period*83/2; Pin <= '1'; wait for clk_period*83/2;
Pin <= '0'; wait for clk_period*84/2; Pin <= '1'; wait for clk_period*84/2;
Pin <= '0'; wait for clk_period*85/2; Pin <= '1'; wait for clk_period*85/2;
Pin <= '0'; wait for clk_period*86/2; Pin <= '1'; wait for clk_period*86/2;
Pin <= '0'; wait for clk_period*87/2; Pin <= '1'; wait for clk_period*87/2;
Pin <= '0'; wait for clk_period*88/2; Pin <= '1'; wait for clk_period*88/2;
Pin <= '0'; wait for clk_period*89/2; Pin <= '1'; wait for clk_period*89/2;
Pin <= '0'; wait for clk_period*90/2; Pin <= '1'; wait for clk_period*90/2;
Pin <= '0'; wait for clk_period*91/2; Pin <= '1'; wait for clk_period*91/2;
Pin <= '0'; wait for clk_period*92/2; Pin <= '1'; wait for clk_period*92/2;
Pin <= '0'; wait for clk_period*93/2; Pin <= '1'; wait for clk_period*93/2;
Pin <= '0'; wait for clk_period*94/2; Pin <= '1'; wait for clk_period*94/2;
Pin <= '0'; wait for clk_period*95/2; Pin <= '1'; wait for clk_period*95/2;
Pin <= '0'; wait for clk_period*96/2; Pin <= '1'; wait for clk_period*96/2;
Pin <= '0'; wait for clk_period*97/2; Pin <= '1'; wait for clk_period*97/2;
Pin <= '0'; wait for clk_period*98/2; Pin <= '1'; wait for clk_period*98/2;
Pin <= '0'; wait for clk_period*99/2; Pin <= '1'; wait for clk_period*99/2;
Pin <= '0'; wait for clk_period*100/2; Pin <= '1'; wait for clk_period*100/2;
Pin <= '0'; wait for clk_period*101/2; Pin <= '1'; wait for clk_period*101/2;
Pin <= '0'; wait for clk_period*102/2; Pin <= '1'; wait for clk_period*102/2;
Pin <= '0'; wait for clk_period*103/2; Pin <= '1'; wait for clk_period*103/2;
Pin <= '0'; wait for clk_period*104/2; Pin <= '1'; wait for clk_period*104/2;
Pin <= '0'; wait for clk_period*105/2; Pin <= '1'; wait for clk_period*105/2;
Pin <= '0'; wait for clk_period*106/2; Pin <= '1'; wait for clk_period*106/2;
Pin <= '0'; wait for clk_period*107/2; Pin <= '1'; wait for clk_period*107/2;
Pin <= '0'; wait for clk_period*108/2; Pin <= '1'; wait for clk_period*108/2;
Pin <= '0'; wait for clk_period*109/2; Pin <= '1'; wait for clk_period*109/2;
Pin <= '0'; wait for clk_period*110/2; Pin <= '1'; wait for clk_period*110/2;
Pin <= '0'; wait for clk_period*111/2; Pin <= '1'; wait for clk_period*111/2;
Pin <= '0'; wait for clk_period*112/2; Pin <= '1'; wait for clk_period*112/2;
Pin <= '0'; wait for clk_period*113/2; Pin <= '1'; wait for clk_period*113/2;
Pin <= '0'; wait for clk_period*114/2; Pin <= '1'; wait for clk_period*114/2;
Pin <= '0'; wait for clk_period*115/2; Pin <= '1'; wait for clk_period*115/2;
Pin <= '0'; wait for clk_period*116/2; Pin <= '1'; wait for clk_period*116/2;
Pin <= '0'; wait for clk_period*117/2; Pin <= '1'; wait for clk_period*117/2;
Pin <= '0'; wait for clk_period*118/2; Pin <= '1'; wait for clk_period*118/2;
Pin <= '0'; wait for clk_period*119/2; Pin <= '1'; wait for clk_period*119/2;
Pin <= '0'; wait for clk_period*120/2; Pin <= '1'; wait for clk_period*120/2;
Pin <= '0'; wait for clk_period*121/2; Pin <= '1'; wait for clk_period*121/2;
Pin <= '0'; wait for clk_period*122/2; Pin <= '1'; wait for clk_period*122/2;
Pin <= '0'; wait for clk_period*123/2; Pin <= '1'; wait for clk_period*123/2;
Pin <= '0'; wait for clk_period*124/2; Pin <= '1'; wait for clk_period*124/2;
Pin <= '0'; wait for clk_period*125/2; Pin <= '1'; wait for clk_period*125/2;
Pin <= '0'; wait for clk_period*126/2; Pin <= '1'; wait for clk_period*126/2;
Pin <= '0'; wait for clk_period*127/2; Pin <= '1'; wait for clk_period*127/2;
Pin <= '0'; wait for clk_period*128/2; Pin <= '1'; wait for clk_period*128/2;
Pin <= '0'; wait for clk_period*129/2; Pin <= '1'; wait for clk_period*129/2;
Pin <= '0'; wait for clk_period*130/2; Pin <= '1'; wait for clk_period*130/2;
Pin <= '0'; wait for clk_period*131/2; Pin <= '1'; wait for clk_period*131/2;
Pin <= '0'; wait for clk_period*132/2; Pin <= '1'; wait for clk_period*132/2;
Pin <= '0'; wait for clk_period*133/2; Pin <= '1'; wait for clk_period*133/2;
Pin <= '0'; wait for clk_period*134/2; Pin <= '1'; wait for clk_period*134/2;
Pin <= '0'; wait for clk_period*135/2; Pin <= '1'; wait for clk_period*135/2;
Pin <= '0'; wait for clk_period*136/2; Pin <= '1'; wait for clk_period*136/2;
Pin <= '0'; wait for clk_period*137/2; Pin <= '1'; wait for clk_period*137/2;
Pin <= '0'; wait for clk_period*138/2; Pin <= '1'; wait for clk_period*138/2;
Pin <= '0'; wait for clk_period*139/2; Pin <= '1'; wait for clk_period*139/2;
Pin <= '0'; wait for clk_period*140/2; Pin <= '1'; wait for clk_period*140/2;
Pin <= '0'; wait for clk_period*141/2; Pin <= '1'; wait for clk_period*141/2;
Pin <= '0'; wait for clk_period*142/2; Pin <= '1'; wait for clk_period*142/2;
Pin <= '0'; wait for clk_period*143/2; Pin <= '1'; wait for clk_period*143/2;
Pin <= '0'; wait for clk_period*144/2; Pin <= '1'; wait for clk_period*144/2;
Pin <= '0'; wait for clk_period*145/2; Pin <= '1'; wait for clk_period*145/2;
Pin <= '0'; wait for clk_period*146/2; Pin <= '1'; wait for clk_period*146/2;
Pin <= '0'; wait for clk_period*147/2; Pin <= '1'; wait for clk_period*147/2;
Pin <= '0'; wait for clk_period*148/2; Pin <= '1'; wait for clk_period*148/2;
Pin <= '0'; wait for clk_period*149/2; Pin <= '1'; wait for clk_period*149/2;
Pin <= '0'; wait for clk_period*150/2; Pin <= '1'; wait for clk_period*150/2;
Pin <= '0'; wait for clk_period*151/2; Pin <= '1'; wait for clk_period*151/2;
Pin <= '0'; wait for clk_period*152/2; Pin <= '1'; wait for clk_period*152/2;
Pin <= '0'; wait for clk_period*153/2; Pin <= '1'; wait for clk_period*153/2;
Pin <= '0'; wait for clk_period*154/2; Pin <= '1'; wait for clk_period*154/2;
Pin <= '0'; wait for clk_period*155/2; Pin <= '1'; wait for clk_period*155/2;
Pin <= '0'; wait for clk_period*156/2; Pin <= '1'; wait for clk_period*156/2;
Pin <= '0'; wait for clk_period*157/2; Pin <= '1'; wait for clk_period*157/2;
Pin <= '0'; wait for clk_period*158/2; Pin <= '1'; wait for clk_period*158/2;
Pin <= '0'; wait for clk_period*159/2; Pin <= '1'; wait for clk_period*159/2;
Pin <= '0'; wait for clk_period*160/2; Pin <= '1'; wait for clk_period*160/2;
Pin <= '0'; wait for clk_period*161/2; Pin <= '1'; wait for clk_period*161/2;
Pin <= '0'; wait for clk_period*162/2; Pin <= '1'; wait for clk_period*162/2;
Pin <= '0'; wait for clk_period*163/2; Pin <= '1'; wait for clk_period*163/2;
Pin <= '0'; wait for clk_period*164/2; Pin <= '1'; wait for clk_period*164/2;
Pin <= '0'; wait for clk_period*165/2; Pin <= '1'; wait for clk_period*165/2;
Pin <= '0'; wait for clk_period*166/2; Pin <= '1'; wait for clk_period*166/2;
Pin <= '0'; wait for clk_period*167/2; Pin <= '1'; wait for clk_period*167/2;
Pin <= '0'; wait for clk_period*168/2; Pin <= '1'; wait for clk_period*168/2;
Pin <= '0'; wait for clk_period*169/2; Pin <= '1'; wait for clk_period*169/2;
Pin <= '0'; wait for clk_period*170/2; Pin <= '1'; wait for clk_period*170/2;
Pin <= '0'; wait for clk_period*171/2; Pin <= '1'; wait for clk_period*171/2;
Pin <= '0'; wait for clk_period*172/2; Pin <= '1'; wait for clk_period*172/2;
Pin <= '0'; wait for clk_period*173/2; Pin <= '1'; wait for clk_period*173/2;
Pin <= '0'; wait for clk_period*174/2; Pin <= '1'; wait for clk_period*174/2;
Pin <= '0'; wait for clk_period*175/2; Pin <= '1'; wait for clk_period*175/2;
Pin <= '0'; wait for clk_period*176/2; Pin <= '1'; wait for clk_period*176/2;
Pin <= '0'; wait for clk_period*177/2; Pin <= '1'; wait for clk_period*177/2;
Pin <= '0'; wait for clk_period*178/2; Pin <= '1'; wait for clk_period*178/2;
Pin <= '0'; wait for clk_period*179/2; Pin <= '1'; wait for clk_period*179/2;
Pin <= '0'; wait for clk_period*180/2; Pin <= '1'; wait for clk_period*180/2;
Pin <= '0'; wait for clk_period*181/2; Pin <= '1'; wait for clk_period*181/2;
Pin <= '0'; wait for clk_period*182/2; Pin <= '1'; wait for clk_period*182/2;
Pin <= '0'; wait for clk_period*183/2; Pin <= '1'; wait for clk_period*183/2;
Pin <= '0'; wait for clk_period*184/2; Pin <= '1'; wait for clk_period*184/2;
Pin <= '0'; wait for clk_period*185/2; Pin <= '1'; wait for clk_period*185/2;
Pin <= '0'; wait for clk_period*186/2; Pin <= '1'; wait for clk_period*186/2;
Pin <= '0'; wait for clk_period*187/2; Pin <= '1'; wait for clk_period*187/2;
Pin <= '0'; wait for clk_period*188/2; Pin <= '1'; wait for clk_period*188/2;
Pin <= '0'; wait for clk_period*189/2; Pin <= '1'; wait for clk_period*189/2;
Pin <= '0'; wait for clk_period*190/2; Pin <= '1'; wait for clk_period*190/2;
Pin <= '0'; wait for clk_period*191/2; Pin <= '1'; wait for clk_period*191/2;
Pin <= '0'; wait for clk_period*192/2; Pin <= '1'; wait for clk_period*192/2;
Pin <= '0'; wait for clk_period*193/2; Pin <= '1'; wait for clk_period*193/2;
Pin <= '0'; wait for clk_period*194/2; Pin <= '1'; wait for clk_period*194/2;
Pin <= '0'; wait for clk_period*195/2; Pin <= '1'; wait for clk_period*195/2;
Pin <= '0'; wait for clk_period*196/2; Pin <= '1'; wait for clk_period*196/2;
Pin <= '0'; wait for clk_period*197/2; Pin <= '1'; wait for clk_period*197/2;
Pin <= '0'; wait for clk_period*198/2; Pin <= '1'; wait for clk_period*198/2;
Pin <= '0'; wait for clk_period*199/2; Pin <= '1'; wait for clk_period*199/2;
Pin <= '0'; wait for clk_period*200/2; Pin <= '1'; wait for clk_period*200/2;
Pin <= '0'; wait for clk_period*201/2; Pin <= '1'; wait for clk_period*201/2;
Pin <= '0'; wait for clk_period*202/2; Pin <= '1'; wait for clk_period*202/2;
Pin <= '0'; wait for clk_period*203/2; Pin <= '1'; wait for clk_period*203/2;
Pin <= '0'; wait for clk_period*204/2; Pin <= '1'; wait for clk_period*204/2;
Pin <= '0'; wait for clk_period*205/2; Pin <= '1'; wait for clk_period*205/2;
Pin <= '0'; wait for clk_period*206/2; Pin <= '1'; wait for clk_period*206/2;
Pin <= '0'; wait for clk_period*207/2; Pin <= '1'; wait for clk_period*207/2;
Pin <= '0'; wait for clk_period*208/2; Pin <= '1'; wait for clk_period*208/2;
Pin <= '0'; wait for clk_period*209/2; Pin <= '1'; wait for clk_period*209/2;
Pin <= '0'; wait for clk_period*210/2; Pin <= '1'; wait for clk_period*210/2;
Pin <= '0'; wait for clk_period*211/2; Pin <= '1'; wait for clk_period*211/2;
Pin <= '0'; wait for clk_period*212/2; Pin <= '1'; wait for clk_period*212/2;
Pin <= '0'; wait for clk_period*213/2; Pin <= '1'; wait for clk_period*213/2;
Pin <= '0'; wait for clk_period*214/2; Pin <= '1'; wait for clk_period*214/2;
Pin <= '0'; wait for clk_period*215/2; Pin <= '1'; wait for clk_period*215/2;
Pin <= '0'; wait for clk_period*216/2; Pin <= '1'; wait for clk_period*216/2;
Pin <= '0'; wait for clk_period*217/2; Pin <= '1'; wait for clk_period*217/2;
Pin <= '0'; wait for clk_period*218/2; Pin <= '1'; wait for clk_period*218/2;
Pin <= '0'; wait for clk_period*219/2; Pin <= '1'; wait for clk_period*219/2;
Pin <= '0'; wait for clk_period*220/2; Pin <= '1'; wait for clk_period*220/2;
Pin <= '0'; wait for clk_period*221/2; Pin <= '1'; wait for clk_period*221/2;
Pin <= '0'; wait for clk_period*222/2; Pin <= '1'; wait for clk_period*222/2;
Pin <= '0'; wait for clk_period*223/2; Pin <= '1'; wait for clk_period*223/2;
Pin <= '0'; wait for clk_period*224/2; Pin <= '1'; wait for clk_period*224/2;
Pin <= '0'; wait for clk_period*225/2; Pin <= '1'; wait for clk_period*225/2;
Pin <= '0'; wait for clk_period*226/2; Pin <= '1'; wait for clk_period*226/2;
Pin <= '0'; wait for clk_period*227/2; Pin <= '1'; wait for clk_period*227/2;
Pin <= '0'; wait for clk_period*228/2; Pin <= '1'; wait for clk_period*228/2;
Pin <= '0'; wait for clk_period*229/2; Pin <= '1'; wait for clk_period*229/2;
Pin <= '0'; wait for clk_period*230/2; Pin <= '1'; wait for clk_period*230/2;
Pin <= '0'; wait for clk_period*231/2; Pin <= '1'; wait for clk_period*231/2;
Pin <= '0'; wait for clk_period*232/2; Pin <= '1'; wait for clk_period*232/2;
Pin <= '0'; wait for clk_period*233/2; Pin <= '1'; wait for clk_period*233/2;
Pin <= '0'; wait for clk_period*234/2; Pin <= '1'; wait for clk_period*234/2;
Pin <= '0'; wait for clk_period*235/2; Pin <= '1'; wait for clk_period*235/2;
Pin <= '0'; wait for clk_period*236/2; Pin <= '1'; wait for clk_period*236/2;
Pin <= '0'; wait for clk_period*237/2; Pin <= '1'; wait for clk_period*237/2;
Pin <= '0'; wait for clk_period*238/2; Pin <= '1'; wait for clk_period*238/2;
Pin <= '0'; wait for clk_period*239/2; Pin <= '1'; wait for clk_period*239/2;
Pin <= '0'; wait for clk_period*240/2; Pin <= '1'; wait for clk_period*240/2;
Pin <= '0'; wait for clk_period*241/2; Pin <= '1'; wait for clk_period*241/2;
Pin <= '0'; wait for clk_period*242/2; Pin <= '1'; wait for clk_period*242/2;
Pin <= '0'; wait for clk_period*243/2; Pin <= '1'; wait for clk_period*243/2;
Pin <= '0'; wait for clk_period*244/2; Pin <= '1'; wait for clk_period*244/2;
Pin <= '0'; wait for clk_period*245/2; Pin <= '1'; wait for clk_period*245/2;
Pin <= '0'; wait for clk_period*246/2; Pin <= '1'; wait for clk_period*246/2;
Pin <= '0'; wait for clk_period*247/2; Pin <= '1'; wait for clk_period*247/2;
Pin <= '0'; wait for clk_period*248/2; Pin <= '1'; wait for clk_period*248/2;
Pin <= '0'; wait for clk_period*249/2; Pin <= '1'; wait for clk_period*249/2;
Pin <= '0'; wait for clk_period*250/2; Pin <= '1'; wait for clk_period*250/2;
Pin <= '0'; wait for clk_period*251/2; Pin <= '1'; wait for clk_period*251/2;
Pin <= '0'; wait for clk_period*252/2; Pin <= '1'; wait for clk_period*252/2;
Pin <= '0'; wait for clk_period*253/2; Pin <= '1'; wait for clk_period*253/2;
Pin <= '0'; wait for clk_period*254/2; Pin <= '1'; wait for clk_period*254/2;
Pin <= '0'; wait for clk_period*255/2; Pin <= '1'; wait for clk_period*255/2;
Pin <= '0'; wait for clk_period*256/2; Pin <= '1'; wait for clk_period*256/2;
Pin <= '0'; wait for clk_period*257/2; Pin <= '1'; wait for clk_period*257/2;
Pin <= '0'; wait for clk_period*258/2; Pin <= '1'; wait for clk_period*258/2;
Pin <= '0'; wait for clk_period*259/2; Pin <= '1'; wait for clk_period*259/2;
Pin <= '0'; wait for clk_period*260/2; Pin <= '1'; wait for clk_period*260/2;
Pin <= '0'; wait for clk_period*261/2; Pin <= '1'; wait for clk_period*261/2;
Pin <= '0'; wait for clk_period*262/2; Pin <= '1'; wait for clk_period*262/2;
Pin <= '0'; wait for clk_period*263/2; Pin <= '1'; wait for clk_period*263/2;
Pin <= '0'; wait for clk_period*264/2; Pin <= '1'; wait for clk_period*264/2;
Pin <= '0'; wait for clk_period*265/2; Pin <= '1'; wait for clk_period*265/2;
Pin <= '0'; wait for clk_period*266/2; Pin <= '1'; wait for clk_period*266/2;
Pin <= '0'; wait for clk_period*267/2; Pin <= '1'; wait for clk_period*267/2;
Pin <= '0'; wait for clk_period*268/2; Pin <= '1'; wait for clk_period*268/2;
Pin <= '0'; wait for clk_period*269/2; Pin <= '1'; wait for clk_period*269/2;
Pin <= '0'; wait for clk_period*270/2; Pin <= '1'; wait for clk_period*270/2;
Pin <= '0'; wait for clk_period*271/2; Pin <= '1'; wait for clk_period*271/2;
Pin <= '0'; wait for clk_period*272/2; Pin <= '1'; wait for clk_period*272/2;
Pin <= '0'; wait for clk_period*273/2; Pin <= '1'; wait for clk_period*273/2;
Pin <= '0'; wait for clk_period*274/2; Pin <= '1'; wait for clk_period*274/2;
Pin <= '0'; wait for clk_period*275/2; Pin <= '1'; wait for clk_period*275/2;
Pin <= '0'; wait for clk_period*276/2; Pin <= '1'; wait for clk_period*276/2;
Pin <= '0'; wait for clk_period*277/2; Pin <= '1'; wait for clk_period*277/2;
Pin <= '0'; wait for clk_period*278/2; Pin <= '1'; wait for clk_period*278/2;
Pin <= '0'; wait for clk_period*279/2; Pin <= '1'; wait for clk_period*279/2;
Pin <= '0'; wait for clk_period*280/2; Pin <= '1'; wait for clk_period*280/2;
Pin <= '0'; wait for clk_period*281/2; Pin <= '1'; wait for clk_period*281/2;
Pin <= '0'; wait for clk_period*282/2; Pin <= '1'; wait for clk_period*282/2;
Pin <= '0'; wait for clk_period*283/2; Pin <= '1'; wait for clk_period*283/2;
Pin <= '0'; wait for clk_period*284/2; Pin <= '1'; wait for clk_period*284/2;
Pin <= '0'; wait for clk_period*285/2; Pin <= '1'; wait for clk_period*285/2;
Pin <= '0'; wait for clk_period*286/2; Pin <= '1'; wait for clk_period*286/2;
Pin <= '0'; wait for clk_period*287/2; Pin <= '1'; wait for clk_period*287/2;
Pin <= '0'; wait for clk_period*288/2; Pin <= '1'; wait for clk_period*288/2;
Pin <= '0'; wait for clk_period*289/2; Pin <= '1'; wait for clk_period*289/2;
Pin <= '0'; wait for clk_period*290/2; Pin <= '1'; wait for clk_period*290/2;
Pin <= '0'; wait for clk_period*291/2; Pin <= '1'; wait for clk_period*291/2;
Pin <= '0'; wait for clk_period*292/2; Pin <= '1'; wait for clk_period*292/2;
Pin <= '0'; wait for clk_period*293/2; Pin <= '1'; wait for clk_period*293/2;
Pin <= '0'; wait for clk_period*294/2; Pin <= '1'; wait for clk_period*294/2;
Pin <= '0'; wait for clk_period*295/2; Pin <= '1'; wait for clk_period*295/2;
Pin <= '0'; wait for clk_period*296/2; Pin <= '1'; wait for clk_period*296/2;
Pin <= '0'; wait for clk_period*297/2; Pin <= '1'; wait for clk_period*297/2;
Pin <= '0'; wait for clk_period*298/2; Pin <= '1'; wait for clk_period*298/2;
Pin <= '0'; wait for clk_period*299/2; Pin <= '1'; wait for clk_period*299/2;
Pin <= '0'; wait for clk_period*300/2; Pin <= '1'; wait for clk_period*300/2;
Pin <= '0'; wait for clk_period*301/2; Pin <= '1'; wait for clk_period*301/2;
Pin <= '0'; wait for clk_period*302/2; Pin <= '1'; wait for clk_period*302/2;
Pin <= '0'; wait for clk_period*303/2; Pin <= '1'; wait for clk_period*303/2;
Pin <= '0'; wait for clk_period*304/2; Pin <= '1'; wait for clk_period*304/2;
Pin <= '0'; wait for clk_period*305/2; Pin <= '1'; wait for clk_period*305/2;
Pin <= '0'; wait for clk_period*306/2; Pin <= '1'; wait for clk_period*306/2;
Pin <= '0'; wait for clk_period*307/2; Pin <= '1'; wait for clk_period*307/2;
Pin <= '0'; wait for clk_period*308/2; Pin <= '1'; wait for clk_period*308/2;
Pin <= '0'; wait for clk_period*309/2; Pin <= '1'; wait for clk_period*309/2;
Pin <= '0'; wait for clk_period*310/2; Pin <= '1'; wait for clk_period*310/2;
Pin <= '0'; wait for clk_period*311/2; Pin <= '1'; wait for clk_period*311/2;
Pin <= '0'; wait for clk_period*312/2; Pin <= '1'; wait for clk_period*312/2;
Pin <= '0'; wait for clk_period*313/2; Pin <= '1'; wait for clk_period*313/2;
Pin <= '0'; wait for clk_period*314/2; Pin <= '1'; wait for clk_period*314/2;
Pin <= '0'; wait for clk_period*315/2; Pin <= '1'; wait for clk_period*315/2;
Pin <= '0'; wait for clk_period*316/2; Pin <= '1'; wait for clk_period*316/2;
Pin <= '0'; wait for clk_period*317/2; Pin <= '1'; wait for clk_period*317/2;
Pin <= '0'; wait for clk_period*318/2; Pin <= '1'; wait for clk_period*318/2;
Pin <= '0'; wait for clk_period*319/2; Pin <= '1'; wait for clk_period*319/2;
Pin <= '0'; wait for clk_period*320/2; Pin <= '1'; wait for clk_period*320/2;
Pin <= '0'; wait for clk_period*321/2; Pin <= '1'; wait for clk_period*321/2;
Pin <= '0'; wait for clk_period*322/2; Pin <= '1'; wait for clk_period*322/2;
Pin <= '0'; wait for clk_period*323/2; Pin <= '1'; wait for clk_period*323/2;
Pin <= '0'; wait for clk_period*324/2; Pin <= '1'; wait for clk_period*324/2;
Pin <= '0'; wait for clk_period*325/2; Pin <= '1'; wait for clk_period*325/2;
Pin <= '0'; wait for clk_period*326/2; Pin <= '1'; wait for clk_period*326/2;
Pin <= '0'; wait for clk_period*327/2; Pin <= '1'; wait for clk_period*327/2;
Pin <= '0'; wait for clk_period*328/2; Pin <= '1'; wait for clk_period*328/2;
Pin <= '0'; wait for clk_period*329/2; Pin <= '1'; wait for clk_period*329/2;
Pin <= '0'; wait for clk_period*330/2; Pin <= '1'; wait for clk_period*330/2;
Pin <= '0'; wait for clk_period*331/2; Pin <= '1'; wait for clk_period*331/2;
Pin <= '0'; wait for clk_period*332/2; Pin <= '1'; wait for clk_period*332/2;
Pin <= '0'; wait for clk_period*333/2; Pin <= '1'; wait for clk_period*333/2;
Pin <= '0'; wait for clk_period*334/2; Pin <= '1'; wait for clk_period*334/2;
Pin <= '0'; wait for clk_period*335/2; Pin <= '1'; wait for clk_period*335/2;
Pin <= '0'; wait for clk_period*336/2; Pin <= '1'; wait for clk_period*336/2;
Pin <= '0'; wait for clk_period*337/2; Pin <= '1'; wait for clk_period*337/2;
Pin <= '0'; wait for clk_period*338/2; Pin <= '1'; wait for clk_period*338/2;
Pin <= '0'; wait for clk_period*339/2; Pin <= '1'; wait for clk_period*339/2;
Pin <= '0'; wait for clk_period*340/2; Pin <= '1'; wait for clk_period*340/2;
Pin <= '0'; wait for clk_period*341/2; Pin <= '1'; wait for clk_period*341/2;
Pin <= '0'; wait for clk_period*342/2; Pin <= '1'; wait for clk_period*342/2;
Pin <= '0'; wait for clk_period*343/2; Pin <= '1'; wait for clk_period*343/2;
Pin <= '0'; wait for clk_period*344/2; Pin <= '1'; wait for clk_period*344/2;
Pin <= '0'; wait for clk_period*345/2; Pin <= '1'; wait for clk_period*345/2;
Pin <= '0'; wait for clk_period*346/2; Pin <= '1'; wait for clk_period*346/2;
Pin <= '0'; wait for clk_period*347/2; Pin <= '1'; wait for clk_period*347/2;
Pin <= '0'; wait for clk_period*348/2; Pin <= '1'; wait for clk_period*348/2;
Pin <= '0'; wait for clk_period*349/2; Pin <= '1'; wait for clk_period*349/2;
Pin <= '0'; wait for clk_period*350/2; Pin <= '1'; wait for clk_period*350/2;
Pin <= '0'; wait for clk_period*351/2; Pin <= '1'; wait for clk_period*351/2;
Pin <= '0'; wait for clk_period*352/2; Pin <= '1'; wait for clk_period*352/2;
Pin <= '0'; wait for clk_period*353/2; Pin <= '1'; wait for clk_period*353/2;
Pin <= '0'; wait for clk_period*354/2; Pin <= '1'; wait for clk_period*354/2;
Pin <= '0'; wait for clk_period*355/2; Pin <= '1'; wait for clk_period*355/2;
Pin <= '0'; wait for clk_period*356/2; Pin <= '1'; wait for clk_period*356/2;
Pin <= '0'; wait for clk_period*357/2; Pin <= '1'; wait for clk_period*357/2;
Pin <= '0'; wait for clk_period*358/2; Pin <= '1'; wait for clk_period*358/2;
Pin <= '0'; wait for clk_period*359/2; Pin <= '1'; wait for clk_period*359/2;
Pin <= '0'; wait for clk_period*360/2; Pin <= '1'; wait for clk_period*360/2;
Pin <= '0'; wait for clk_period*361/2; Pin <= '1'; wait for clk_period*361/2;
Pin <= '0'; wait for clk_period*362/2; Pin <= '1'; wait for clk_period*362/2;
Pin <= '0'; wait for clk_period*363/2; Pin <= '1'; wait for clk_period*363/2;
Pin <= '0'; wait for clk_period*364/2; Pin <= '1'; wait for clk_period*364/2;
Pin <= '0'; wait for clk_period*365/2; Pin <= '1'; wait for clk_period*365/2;
Pin <= '0'; wait for clk_period*366/2; Pin <= '1'; wait for clk_period*366/2;
Pin <= '0'; wait for clk_period*367/2; Pin <= '1'; wait for clk_period*367/2;
Pin <= '0'; wait for clk_period*368/2; Pin <= '1'; wait for clk_period*368/2;
Pin <= '0'; wait for clk_period*369/2; Pin <= '1'; wait for clk_period*369/2;
Pin <= '0'; wait for clk_period*370/2; Pin <= '1'; wait for clk_period*370/2;
Pin <= '0'; wait for clk_period*371/2; Pin <= '1'; wait for clk_period*371/2;
Pin <= '0'; wait for clk_period*372/2; Pin <= '1'; wait for clk_period*372/2;
Pin <= '0'; wait for clk_period*373/2; Pin <= '1'; wait for clk_period*373/2;
Pin <= '0'; wait for clk_period*374/2; Pin <= '1'; wait for clk_period*374/2;
Pin <= '0'; wait for clk_period*375/2; Pin <= '1'; wait for clk_period*375/2;
Pin <= '0'; wait for clk_period*376/2; Pin <= '1'; wait for clk_period*376/2;
Pin <= '0'; wait for clk_period*377/2; Pin <= '1'; wait for clk_period*377/2;
Pin <= '0'; wait for clk_period*378/2; Pin <= '1'; wait for clk_period*378/2;
Pin <= '0'; wait for clk_period*379/2; Pin <= '1'; wait for clk_period*379/2;
Pin <= '0'; wait for clk_period*380/2; Pin <= '1'; wait for clk_period*380/2;
Pin <= '0'; wait for clk_period*381/2; Pin <= '1'; wait for clk_period*381/2;
Pin <= '0'; wait for clk_period*382/2; Pin <= '1'; wait for clk_period*382/2;
Pin <= '0'; wait for clk_period*383/2; Pin <= '1'; wait for clk_period*383/2;
Pin <= '0'; wait for clk_period*384/2; Pin <= '1'; wait for clk_period*384/2;
Pin <= '0'; wait for clk_period*385/2; Pin <= '1'; wait for clk_period*385/2;
Pin <= '0'; wait for clk_period*386/2; Pin <= '1'; wait for clk_period*386/2;
Pin <= '0'; wait for clk_period*387/2; Pin <= '1'; wait for clk_period*387/2;
Pin <= '0'; wait for clk_period*388/2; Pin <= '1'; wait for clk_period*388/2;
Pin <= '0'; wait for clk_period*389/2; Pin <= '1'; wait for clk_period*389/2;
Pin <= '0'; wait for clk_period*390/2; Pin <= '1'; wait for clk_period*390/2;
Pin <= '0'; wait for clk_period*391/2; Pin <= '1'; wait for clk_period*391/2;
Pin <= '0'; wait for clk_period*392/2; Pin <= '1'; wait for clk_period*392/2;
Pin <= '0'; wait for clk_period*393/2; Pin <= '1'; wait for clk_period*393/2;
Pin <= '0'; wait for clk_period*394/2; Pin <= '1'; wait for clk_period*394/2;
Pin <= '0'; wait for clk_period*395/2; Pin <= '1'; wait for clk_period*395/2;
Pin <= '0'; wait for clk_period*396/2; Pin <= '1'; wait for clk_period*396/2;
Pin <= '0'; wait for clk_period*397/2; Pin <= '1'; wait for clk_period*397/2;
Pin <= '0'; wait for clk_period*398/2; Pin <= '1'; wait for clk_period*398/2;
Pin <= '0'; wait for clk_period*399/2; Pin <= '1'; wait for clk_period*399/2;
Pin <= '0'; wait for clk_period*400/2; Pin <= '1'; wait for clk_period*400/2;
Pin <= '0'; wait for clk_period*401/2; Pin <= '1'; wait for clk_period*401/2;
Pin <= '0'; wait for clk_period*402/2; Pin <= '1'; wait for clk_period*402/2;
Pin <= '0'; wait for clk_period*403/2; Pin <= '1'; wait for clk_period*403/2;
Pin <= '0'; wait for clk_period*404/2; Pin <= '1'; wait for clk_period*404/2;
Pin <= '0'; wait for clk_period*405/2; Pin <= '1'; wait for clk_period*405/2;
Pin <= '0'; wait for clk_period*406/2; Pin <= '1'; wait for clk_period*406/2;
Pin <= '0'; wait for clk_period*407/2; Pin <= '1'; wait for clk_period*407/2;
Pin <= '0'; wait for clk_period*408/2; Pin <= '1'; wait for clk_period*408/2;
Pin <= '0'; wait for clk_period*409/2; Pin <= '1'; wait for clk_period*409/2;
Pin <= '0'; wait for clk_period*410/2; Pin <= '1'; wait for clk_period*410/2;
Pin <= '0'; wait for clk_period*411/2; Pin <= '1'; wait for clk_period*411/2;
Pin <= '0'; wait for clk_period*412/2; Pin <= '1'; wait for clk_period*412/2;
Pin <= '0'; wait for clk_period*413/2; Pin <= '1'; wait for clk_period*413/2;
Pin <= '0'; wait for clk_period*414/2; Pin <= '1'; wait for clk_period*414/2;
Pin <= '0'; wait for clk_period*415/2; Pin <= '1'; wait for clk_period*415/2;
Pin <= '0'; wait for clk_period*416/2; Pin <= '1'; wait for clk_period*416/2;
Pin <= '0'; wait for clk_period*417/2; Pin <= '1'; wait for clk_period*417/2;
Pin <= '0'; wait for clk_period*418/2; Pin <= '1'; wait for clk_period*418/2;
Pin <= '0'; wait for clk_period*419/2; Pin <= '1'; wait for clk_period*419/2;
Pin <= '0'; wait for clk_period*420/2; Pin <= '1'; wait for clk_period*420/2;
Pin <= '0'; wait for clk_period*421/2; Pin <= '1'; wait for clk_period*421/2;
Pin <= '0'; wait for clk_period*422/2; Pin <= '1'; wait for clk_period*422/2;
Pin <= '0'; wait for clk_period*423/2; Pin <= '1'; wait for clk_period*423/2;
Pin <= '0'; wait for clk_period*424/2; Pin <= '1'; wait for clk_period*424/2;
Pin <= '0'; wait for clk_period*425/2; Pin <= '1'; wait for clk_period*425/2;
Pin <= '0'; wait for clk_period*426/2; Pin <= '1'; wait for clk_period*426/2;
Pin <= '0'; wait for clk_period*427/2; Pin <= '1'; wait for clk_period*427/2;
Pin <= '0'; wait for clk_period*428/2; Pin <= '1'; wait for clk_period*428/2;
Pin <= '0'; wait for clk_period*429/2; Pin <= '1'; wait for clk_period*429/2;
Pin <= '0'; wait for clk_period*430/2; Pin <= '1'; wait for clk_period*430/2;
Pin <= '0'; wait for clk_period*431/2; Pin <= '1'; wait for clk_period*431/2;
Pin <= '0'; wait for clk_period*432/2; Pin <= '1'; wait for clk_period*432/2;
Pin <= '0'; wait for clk_period*433/2; Pin <= '1'; wait for clk_period*433/2;
Pin <= '0'; wait for clk_period*434/2; Pin <= '1'; wait for clk_period*434/2;
Pin <= '0'; wait for clk_period*435/2; Pin <= '1'; wait for clk_period*435/2;
Pin <= '0'; wait for clk_period*436/2; Pin <= '1'; wait for clk_period*436/2;
Pin <= '0'; wait for clk_period*437/2; Pin <= '1'; wait for clk_period*437/2;
Pin <= '0'; wait for clk_period*438/2; Pin <= '1'; wait for clk_period*438/2;
Pin <= '0'; wait for clk_period*439/2; Pin <= '1'; wait for clk_period*439/2;
Pin <= '0'; wait for clk_period*440/2; Pin <= '1'; wait for clk_period*440/2;
Pin <= '0'; wait for clk_period*441/2; Pin <= '1'; wait for clk_period*441/2;
Pin <= '0'; wait for clk_period*442/2; Pin <= '1'; wait for clk_period*442/2;
Pin <= '0'; wait for clk_period*443/2; Pin <= '1'; wait for clk_period*443/2;
Pin <= '0'; wait for clk_period*444/2; Pin <= '1'; wait for clk_period*444/2;
Pin <= '0'; wait for clk_period*445/2; Pin <= '1'; wait for clk_period*445/2;
Pin <= '0'; wait for clk_period*446/2; Pin <= '1'; wait for clk_period*446/2;
Pin <= '0'; wait for clk_period*447/2; Pin <= '1'; wait for clk_period*447/2;
Pin <= '0'; wait for clk_period*448/2; Pin <= '1'; wait for clk_period*448/2;
Pin <= '0'; wait for clk_period*449/2; Pin <= '1'; wait for clk_period*449/2;
Pin <= '0'; wait for clk_period*450/2; Pin <= '1'; wait for clk_period*450/2;
Pin <= '0'; wait for clk_period*451/2; Pin <= '1'; wait for clk_period*451/2;
Pin <= '0'; wait for clk_period*452/2; Pin <= '1'; wait for clk_period*452/2;
Pin <= '0'; wait for clk_period*453/2; Pin <= '1'; wait for clk_period*453/2;
Pin <= '0'; wait for clk_period*454/2; Pin <= '1'; wait for clk_period*454/2;
Pin <= '0'; wait for clk_period*455/2; Pin <= '1'; wait for clk_period*455/2;
Pin <= '0'; wait for clk_period*456/2; Pin <= '1'; wait for clk_period*456/2;
Pin <= '0'; wait for clk_period*457/2; Pin <= '1'; wait for clk_period*457/2;
Pin <= '0'; wait for clk_period*458/2; Pin <= '1'; wait for clk_period*458/2;
Pin <= '0'; wait for clk_period*459/2; Pin <= '1'; wait for clk_period*459/2;
Pin <= '0'; wait for clk_period*460/2; Pin <= '1'; wait for clk_period*460/2;
Pin <= '0'; wait for clk_period*461/2; Pin <= '1'; wait for clk_period*461/2;
Pin <= '0'; wait for clk_period*462/2; Pin <= '1'; wait for clk_period*462/2;
Pin <= '0'; wait for clk_period*463/2; Pin <= '1'; wait for clk_period*463/2;
Pin <= '0'; wait for clk_period*464/2; Pin <= '1'; wait for clk_period*464/2;
Pin <= '0'; wait for clk_period*465/2; Pin <= '1'; wait for clk_period*465/2;
Pin <= '0'; wait for clk_period*466/2; Pin <= '1'; wait for clk_period*466/2;
Pin <= '0'; wait for clk_period*467/2; Pin <= '1'; wait for clk_period*467/2;
Pin <= '0'; wait for clk_period*468/2; Pin <= '1'; wait for clk_period*468/2;
Pin <= '0'; wait for clk_period*469/2; Pin <= '1'; wait for clk_period*469/2;
Pin <= '0'; wait for clk_period*470/2; Pin <= '1'; wait for clk_period*470/2;
Pin <= '0'; wait for clk_period*471/2; Pin <= '1'; wait for clk_period*471/2;
Pin <= '0'; wait for clk_period*472/2; Pin <= '1'; wait for clk_period*472/2;
Pin <= '0'; wait for clk_period*473/2; Pin <= '1'; wait for clk_period*473/2;
Pin <= '0'; wait for clk_period*474/2; Pin <= '1'; wait for clk_period*474/2;
Pin <= '0'; wait for clk_period*475/2; Pin <= '1'; wait for clk_period*475/2;
Pin <= '0'; wait for clk_period*476/2; Pin <= '1'; wait for clk_period*476/2;
Pin <= '0'; wait for clk_period*477/2; Pin <= '1'; wait for clk_period*477/2;
Pin <= '0'; wait for clk_period*478/2; Pin <= '1'; wait for clk_period*478/2;
Pin <= '0'; wait for clk_period*479/2; Pin <= '1'; wait for clk_period*479/2;
Pin <= '0'; wait for clk_period*480/2; Pin <= '1'; wait for clk_period*480/2;
Pin <= '0'; wait for clk_period*481/2; Pin <= '1'; wait for clk_period*481/2;
Pin <= '0'; wait for clk_period*482/2; Pin <= '1'; wait for clk_period*482/2;
Pin <= '0'; wait for clk_period*483/2; Pin <= '1'; wait for clk_period*483/2;
Pin <= '0'; wait for clk_period*484/2; Pin <= '1'; wait for clk_period*484/2;
Pin <= '0'; wait for clk_period*485/2; Pin <= '1'; wait for clk_period*485/2;
Pin <= '0'; wait for clk_period*486/2; Pin <= '1'; wait for clk_period*486/2;
Pin <= '0'; wait for clk_period*487/2; Pin <= '1'; wait for clk_period*487/2;
Pin <= '0'; wait for clk_period*488/2; Pin <= '1'; wait for clk_period*488/2;
Pin <= '0'; wait for clk_period*489/2; Pin <= '1'; wait for clk_period*489/2;
Pin <= '0'; wait for clk_period*490/2; Pin <= '1'; wait for clk_period*490/2;
Pin <= '0'; wait for clk_period*491/2; Pin <= '1'; wait for clk_period*491/2;
Pin <= '0'; wait for clk_period*492/2; Pin <= '1'; wait for clk_period*492/2;
Pin <= '0'; wait for clk_period*493/2; Pin <= '1'; wait for clk_period*493/2;
Pin <= '0'; wait for clk_period*494/2; Pin <= '1'; wait for clk_period*494/2;
Pin <= '0'; wait for clk_period*495/2; Pin <= '1'; wait for clk_period*495/2;
Pin <= '0'; wait for clk_period*496/2; Pin <= '1'; wait for clk_period*496/2;
Pin <= '0'; wait for clk_period*497/2; Pin <= '1'; wait for clk_period*497/2;
Pin <= '0'; wait for clk_period*498/2; Pin <= '1'; wait for clk_period*498/2;
Pin <= '0'; wait for clk_period*499/2; Pin <= '1'; wait for clk_period*499/2;
Pin <= '0'; wait for clk_period*500/2; Pin <= '1'; wait for clk_period*500/2;
Pin <= '0'; wait for clk_period*501/2; Pin <= '1'; wait for clk_period*501/2;
Pin <= '0'; wait for clk_period*502/2; Pin <= '1'; wait for clk_period*502/2;
Pin <= '0'; wait for clk_period*503/2; Pin <= '1'; wait for clk_period*503/2;
Pin <= '0'; wait for clk_period*504/2; Pin <= '1'; wait for clk_period*504/2;
Pin <= '0'; wait for clk_period*505/2; Pin <= '1'; wait for clk_period*505/2;
Pin <= '0'; wait for clk_period*506/2; Pin <= '1'; wait for clk_period*506/2;
Pin <= '0'; wait for clk_period*507/2; Pin <= '1'; wait for clk_period*507/2;
Pin <= '0'; wait for clk_period*508/2; Pin <= '1'; wait for clk_period*508/2;
Pin <= '0'; wait for clk_period*509/2; Pin <= '1'; wait for clk_period*509/2;
Pin <= '0'; wait for clk_period*510/2; Pin <= '1'; wait for clk_period*510/2;
Pin <= '0'; wait for clk_period*511/2; Pin <= '1'; wait for clk_period*511/2;
Pin <= '0'; wait for clk_period*512/2; Pin <= '1'; wait for clk_period*512/2;
Pin <= '0'; wait for clk_period*513/2; Pin <= '1'; wait for clk_period*513/2;
Pin <= '0'; wait for clk_period*514/2; Pin <= '1'; wait for clk_period*514/2;
Pin <= '0'; wait for clk_period*515/2; Pin <= '1'; wait for clk_period*515/2;
Pin <= '0'; wait for clk_period*516/2; Pin <= '1'; wait for clk_period*516/2;
Pin <= '0'; wait for clk_period*517/2; Pin <= '1'; wait for clk_period*517/2;
Pin <= '0'; wait for clk_period*518/2; Pin <= '1'; wait for clk_period*518/2;
Pin <= '0'; wait for clk_period*519/2; Pin <= '1'; wait for clk_period*519/2;
Pin <= '0'; wait for clk_period*520/2; Pin <= '1'; wait for clk_period*520/2;
Pin <= '0'; wait for clk_period*521/2; Pin <= '1'; wait for clk_period*521/2;
Pin <= '0'; wait for clk_period*522/2; Pin <= '1'; wait for clk_period*522/2;
Pin <= '0'; wait for clk_period*523/2; Pin <= '1'; wait for clk_period*523/2;
Pin <= '0'; wait for clk_period*524/2; Pin <= '1'; wait for clk_period*524/2;
Pin <= '0'; wait for clk_period*525/2; Pin <= '1'; wait for clk_period*525/2;
Pin <= '0'; wait for clk_period*526/2; Pin <= '1'; wait for clk_period*526/2;
Pin <= '0'; wait for clk_period*527/2; Pin <= '1'; wait for clk_period*527/2;
Pin <= '0'; wait for clk_period*528/2; Pin <= '1'; wait for clk_period*528/2;
Pin <= '0'; wait for clk_period*529/2; Pin <= '1'; wait for clk_period*529/2;
Pin <= '0'; wait for clk_period*530/2; Pin <= '1'; wait for clk_period*530/2;
Pin <= '0'; wait for clk_period*531/2; Pin <= '1'; wait for clk_period*531/2;
Pin <= '0'; wait for clk_period*532/2; Pin <= '1'; wait for clk_period*532/2;
Pin <= '0'; wait for clk_period*533/2; Pin <= '1'; wait for clk_period*533/2;
Pin <= '0'; wait for clk_period*534/2; Pin <= '1'; wait for clk_period*534/2;
Pin <= '0'; wait for clk_period*535/2; Pin <= '1'; wait for clk_period*535/2;
Pin <= '0'; wait for clk_period*536/2; Pin <= '1'; wait for clk_period*536/2;
Pin <= '0'; wait for clk_period*537/2; Pin <= '1'; wait for clk_period*537/2;
Pin <= '0'; wait for clk_period*538/2; Pin <= '1'; wait for clk_period*538/2;
Pin <= '0'; wait for clk_period*539/2; Pin <= '1'; wait for clk_period*539/2;
Pin <= '0'; wait for clk_period*540/2; Pin <= '1'; wait for clk_period*540/2;
Pin <= '0'; wait for clk_period*541/2; Pin <= '1'; wait for clk_period*541/2;
Pin <= '0'; wait for clk_period*542/2; Pin <= '1'; wait for clk_period*542/2;
Pin <= '0'; wait for clk_period*543/2; Pin <= '1'; wait for clk_period*543/2;
Pin <= '0'; wait for clk_period*544/2; Pin <= '1'; wait for clk_period*544/2;
Pin <= '0'; wait for clk_period*545/2; Pin <= '1'; wait for clk_period*545/2;
Pin <= '0'; wait for clk_period*546/2; Pin <= '1'; wait for clk_period*546/2;
Pin <= '0'; wait for clk_period*547/2; Pin <= '1'; wait for clk_period*547/2;
Pin <= '0'; wait for clk_period*548/2; Pin <= '1'; wait for clk_period*548/2;
Pin <= '0'; wait for clk_period*549/2; Pin <= '1'; wait for clk_period*549/2;
Pin <= '0'; wait for clk_period*550/2; Pin <= '1'; wait for clk_period*550/2;
Pin <= '0'; wait for clk_period*551/2; Pin <= '1'; wait for clk_period*551/2;
Pin <= '0'; wait for clk_period*552/2; Pin <= '1'; wait for clk_period*552/2;
Pin <= '0'; wait for clk_period*553/2; Pin <= '1'; wait for clk_period*553/2;
Pin <= '0'; wait for clk_period*554/2; Pin <= '1'; wait for clk_period*554/2;
Pin <= '0'; wait for clk_period*555/2; Pin <= '1'; wait for clk_period*555/2;
Pin <= '0'; wait for clk_period*556/2; Pin <= '1'; wait for clk_period*556/2;
Pin <= '0'; wait for clk_period*557/2; Pin <= '1'; wait for clk_period*557/2;
Pin <= '0'; wait for clk_period*558/2; Pin <= '1'; wait for clk_period*558/2;
Pin <= '0'; wait for clk_period*559/2; Pin <= '1'; wait for clk_period*559/2;
Pin <= '0'; wait for clk_period*560/2; Pin <= '1'; wait for clk_period*560/2;
Pin <= '0'; wait for clk_period*561/2; Pin <= '1'; wait for clk_period*561/2;
Pin <= '0'; wait for clk_period*562/2; Pin <= '1'; wait for clk_period*562/2;
Pin <= '0'; wait for clk_period*563/2; Pin <= '1'; wait for clk_period*563/2;
Pin <= '0'; wait for clk_period*564/2; Pin <= '1'; wait for clk_period*564/2;
Pin <= '0'; wait for clk_period*565/2; Pin <= '1'; wait for clk_period*565/2;
Pin <= '0'; wait for clk_period*566/2; Pin <= '1'; wait for clk_period*566/2;
Pin <= '0'; wait for clk_period*567/2; Pin <= '1'; wait for clk_period*567/2;
Pin <= '0'; wait for clk_period*568/2; Pin <= '1'; wait for clk_period*568/2;
Pin <= '0'; wait for clk_period*569/2; Pin <= '1'; wait for clk_period*569/2;
Pin <= '0'; wait for clk_period*570/2; Pin <= '1'; wait for clk_period*570/2;
Pin <= '0'; wait for clk_period*571/2; Pin <= '1'; wait for clk_period*571/2;
Pin <= '0'; wait for clk_period*572/2; Pin <= '1'; wait for clk_period*572/2;
Pin <= '0'; wait for clk_period*573/2; Pin <= '1'; wait for clk_period*573/2;
Pin <= '0'; wait for clk_period*574/2; Pin <= '1'; wait for clk_period*574/2;
Pin <= '0'; wait for clk_period*575/2; Pin <= '1'; wait for clk_period*575/2;
Pin <= '0'; wait for clk_period*576/2; Pin <= '1'; wait for clk_period*576/2;
Pin <= '0'; wait for clk_period*577/2; Pin <= '1'; wait for clk_period*577/2;
Pin <= '0'; wait for clk_period*578/2; Pin <= '1'; wait for clk_period*578/2;
Pin <= '0'; wait for clk_period*579/2; Pin <= '1'; wait for clk_period*579/2;
Pin <= '0'; wait for clk_period*580/2; Pin <= '1'; wait for clk_period*580/2;
Pin <= '0'; wait for clk_period*581/2; Pin <= '1'; wait for clk_period*581/2;
Pin <= '0'; wait for clk_period*582/2; Pin <= '1'; wait for clk_period*582/2;
Pin <= '0'; wait for clk_period*583/2; Pin <= '1'; wait for clk_period*583/2;
Pin <= '0'; wait for clk_period*584/2; Pin <= '1'; wait for clk_period*584/2;
Pin <= '0'; wait for clk_period*585/2; Pin <= '1'; wait for clk_period*585/2;
Pin <= '0'; wait for clk_period*586/2; Pin <= '1'; wait for clk_period*586/2;
Pin <= '0'; wait for clk_period*587/2; Pin <= '1'; wait for clk_period*587/2;
Pin <= '0'; wait for clk_period*588/2; Pin <= '1'; wait for clk_period*588/2;
Pin <= '0'; wait for clk_period*589/2; Pin <= '1'; wait for clk_period*589/2;
Pin <= '0'; wait for clk_period*590/2; Pin <= '1'; wait for clk_period*590/2;
Pin <= '0'; wait for clk_period*591/2; Pin <= '1'; wait for clk_period*591/2;
Pin <= '0'; wait for clk_period*592/2; Pin <= '1'; wait for clk_period*592/2;
Pin <= '0'; wait for clk_period*593/2; Pin <= '1'; wait for clk_period*593/2;
Pin <= '0'; wait for clk_period*594/2; Pin <= '1'; wait for clk_period*594/2;
Pin <= '0'; wait for clk_period*595/2; Pin <= '1'; wait for clk_period*595/2;
Pin <= '0'; wait for clk_period*596/2; Pin <= '1'; wait for clk_period*596/2;
Pin <= '0'; wait for clk_period*597/2; Pin <= '1'; wait for clk_period*597/2;
Pin <= '0'; wait for clk_period*598/2; Pin <= '1'; wait for clk_period*598/2;
Pin <= '0'; wait for clk_period*599/2; Pin <= '1'; wait for clk_period*599/2;
Pin <= '0'; wait for clk_period*600/2; Pin <= '1'; wait for clk_period*600/2;
Pin <= '0'; wait for clk_period*601/2; Pin <= '1'; wait for clk_period*601/2;
Pin <= '0'; wait for clk_period*602/2; Pin <= '1'; wait for clk_period*602/2;
Pin <= '0'; wait for clk_period*603/2; Pin <= '1'; wait for clk_period*603/2;
Pin <= '0'; wait for clk_period*604/2; Pin <= '1'; wait for clk_period*604/2;
Pin <= '0'; wait for clk_period*605/2; Pin <= '1'; wait for clk_period*605/2;
Pin <= '0'; wait for clk_period*606/2; Pin <= '1'; wait for clk_period*606/2;
Pin <= '0'; wait for clk_period*607/2; Pin <= '1'; wait for clk_period*607/2;
Pin <= '0'; wait for clk_period*608/2; Pin <= '1'; wait for clk_period*608/2;
Pin <= '0'; wait for clk_period*609/2; Pin <= '1'; wait for clk_period*609/2;
Pin <= '0'; wait for clk_period*610/2; Pin <= '1'; wait for clk_period*610/2;
Pin <= '0'; wait for clk_period*611/2; Pin <= '1'; wait for clk_period*611/2;
Pin <= '0'; wait for clk_period*612/2; Pin <= '1'; wait for clk_period*612/2;
Pin <= '0'; wait for clk_period*613/2; Pin <= '1'; wait for clk_period*613/2;
Pin <= '0'; wait for clk_period*614/2; Pin <= '1'; wait for clk_period*614/2;
Pin <= '0'; wait for clk_period*615/2; Pin <= '1'; wait for clk_period*615/2;
Pin <= '0'; wait for clk_period*616/2; Pin <= '1'; wait for clk_period*616/2;
Pin <= '0'; wait for clk_period*617/2; Pin <= '1'; wait for clk_period*617/2;
Pin <= '0'; wait for clk_period*618/2; Pin <= '1'; wait for clk_period*618/2;
Pin <= '0'; wait for clk_period*619/2; Pin <= '1'; wait for clk_period*619/2;
Pin <= '0'; wait for clk_period*620/2; Pin <= '1'; wait for clk_period*620/2;
Pin <= '0'; wait for clk_period*621/2; Pin <= '1'; wait for clk_period*621/2;
Pin <= '0'; wait for clk_period*622/2; Pin <= '1'; wait for clk_period*622/2;
Pin <= '0'; wait for clk_period*623/2; Pin <= '1'; wait for clk_period*623/2;
Pin <= '0'; wait for clk_period*624/2; Pin <= '1'; wait for clk_period*624/2;
Pin <= '0'; wait for clk_period*625/2; Pin <= '1'; wait for clk_period*625/2;
Pin <= '0'; wait for clk_period*626/2; Pin <= '1'; wait for clk_period*626/2;
Pin <= '0'; wait for clk_period*627/2; Pin <= '1'; wait for clk_period*627/2;
Pin <= '0'; wait for clk_period*628/2; Pin <= '1'; wait for clk_period*628/2;
Pin <= '0'; wait for clk_period*629/2; Pin <= '1'; wait for clk_period*629/2;
Pin <= '0'; wait for clk_period*630/2; Pin <= '1'; wait for clk_period*630/2;
Pin <= '0'; wait for clk_period*631/2; Pin <= '1'; wait for clk_period*631/2;
Pin <= '0'; wait for clk_period*632/2; Pin <= '1'; wait for clk_period*632/2;
Pin <= '0'; wait for clk_period*633/2; Pin <= '1'; wait for clk_period*633/2;
Pin <= '0'; wait for clk_period*634/2; Pin <= '1'; wait for clk_period*634/2;
Pin <= '0'; wait for clk_period*635/2; Pin <= '1'; wait for clk_period*635/2;
Pin <= '0'; wait for clk_period*636/2; Pin <= '1'; wait for clk_period*636/2;
Pin <= '0'; wait for clk_period*637/2; Pin <= '1'; wait for clk_period*637/2;
Pin <= '0'; wait for clk_period*638/2; Pin <= '1'; wait for clk_period*638/2;
Pin <= '0'; wait for clk_period*639/2; Pin <= '1'; wait for clk_period*639/2;
Pin <= '0'; wait for clk_period*640/2; Pin <= '1'; wait for clk_period*640/2;
Pin <= '0'; wait for clk_period*641/2; Pin <= '1'; wait for clk_period*641/2;
Pin <= '0'; wait for clk_period*642/2; Pin <= '1'; wait for clk_period*642/2;
Pin <= '0'; wait for clk_period*643/2; Pin <= '1'; wait for clk_period*643/2;
Pin <= '0'; wait for clk_period*644/2; Pin <= '1'; wait for clk_period*644/2;
Pin <= '0'; wait for clk_period*645/2; Pin <= '1'; wait for clk_period*645/2;
Pin <= '0'; wait for clk_period*646/2; Pin <= '1'; wait for clk_period*646/2;
Pin <= '0'; wait for clk_period*647/2; Pin <= '1'; wait for clk_period*647/2;
Pin <= '0'; wait for clk_period*648/2; Pin <= '1'; wait for clk_period*648/2;
Pin <= '0'; wait for clk_period*649/2; Pin <= '1'; wait for clk_period*649/2;
Pin <= '0'; wait for clk_period*650/2; Pin <= '1'; wait for clk_period*650/2;
Pin <= '0'; wait for clk_period*651/2; Pin <= '1'; wait for clk_period*651/2;
Pin <= '0'; wait for clk_period*652/2; Pin <= '1'; wait for clk_period*652/2;
Pin <= '0'; wait for clk_period*653/2; Pin <= '1'; wait for clk_period*653/2;
Pin <= '0'; wait for clk_period*654/2; Pin <= '1'; wait for clk_period*654/2;
Pin <= '0'; wait for clk_period*655/2; Pin <= '1'; wait for clk_period*655/2;
Pin <= '0'; wait for clk_period*656/2; Pin <= '1'; wait for clk_period*656/2;
Pin <= '0'; wait for clk_period*657/2; Pin <= '1'; wait for clk_period*657/2;
Pin <= '0'; wait for clk_period*658/2; Pin <= '1'; wait for clk_period*658/2;
Pin <= '0'; wait for clk_period*659/2; Pin <= '1'; wait for clk_period*659/2;
Pin <= '0'; wait for clk_period*660/2; Pin <= '1'; wait for clk_period*660/2;
Pin <= '0'; wait for clk_period*661/2; Pin <= '1'; wait for clk_period*661/2;
Pin <= '0'; wait for clk_period*662/2; Pin <= '1'; wait for clk_period*662/2;
Pin <= '0'; wait for clk_period*663/2; Pin <= '1'; wait for clk_period*663/2;
Pin <= '0'; wait for clk_period*664/2; Pin <= '1'; wait for clk_period*664/2;
Pin <= '0'; wait for clk_period*665/2; Pin <= '1'; wait for clk_period*665/2;
Pin <= '0'; wait for clk_period*666/2; Pin <= '1'; wait for clk_period*666/2;
Pin <= '0'; wait for clk_period*667/2; Pin <= '1'; wait for clk_period*667/2;
Pin <= '0'; wait for clk_period*668/2; Pin <= '1'; wait for clk_period*668/2;
Pin <= '0'; wait for clk_period*669/2; Pin <= '1'; wait for clk_period*669/2;
Pin <= '0'; wait for clk_period*670/2; Pin <= '1'; wait for clk_period*670/2;
Pin <= '0'; wait for clk_period*671/2; Pin <= '1'; wait for clk_period*671/2;
Pin <= '0'; wait for clk_period*672/2; Pin <= '1'; wait for clk_period*672/2;
Pin <= '0'; wait for clk_period*673/2; Pin <= '1'; wait for clk_period*673/2;
Pin <= '0'; wait for clk_period*674/2; Pin <= '1'; wait for clk_period*674/2;
Pin <= '0'; wait for clk_period*675/2; Pin <= '1'; wait for clk_period*675/2;
Pin <= '0'; wait for clk_period*676/2; Pin <= '1'; wait for clk_period*676/2;
Pin <= '0'; wait for clk_period*677/2; Pin <= '1'; wait for clk_period*677/2;
Pin <= '0'; wait for clk_period*678/2; Pin <= '1'; wait for clk_period*678/2;
Pin <= '0'; wait for clk_period*679/2; Pin <= '1'; wait for clk_period*679/2;
Pin <= '0'; wait for clk_period*680/2; Pin <= '1'; wait for clk_period*680/2;
Pin <= '0'; wait for clk_period*681/2; Pin <= '1'; wait for clk_period*681/2;
Pin <= '0'; wait for clk_period*682/2; Pin <= '1'; wait for clk_period*682/2;
Pin <= '0'; wait for clk_period*683/2; Pin <= '1'; wait for clk_period*683/2;
Pin <= '0'; wait for clk_period*684/2; Pin <= '1'; wait for clk_period*684/2;
Pin <= '0'; wait for clk_period*685/2; Pin <= '1'; wait for clk_period*685/2;
Pin <= '0'; wait for clk_period*686/2; Pin <= '1'; wait for clk_period*686/2;
Pin <= '0'; wait for clk_period*687/2; Pin <= '1'; wait for clk_period*687/2;
Pin <= '0'; wait for clk_period*688/2; Pin <= '1'; wait for clk_period*688/2;
Pin <= '0'; wait for clk_period*689/2; Pin <= '1'; wait for clk_period*689/2;
Pin <= '0'; wait for clk_period*690/2; Pin <= '1'; wait for clk_period*690/2;
Pin <= '0'; wait for clk_period*691/2; Pin <= '1'; wait for clk_period*691/2;
Pin <= '0'; wait for clk_period*692/2; Pin <= '1'; wait for clk_period*692/2;
Pin <= '0'; wait for clk_period*693/2; Pin <= '1'; wait for clk_period*693/2;
Pin <= '0'; wait for clk_period*694/2; Pin <= '1'; wait for clk_period*694/2;
Pin <= '0'; wait for clk_period*695/2; Pin <= '1'; wait for clk_period*695/2;
Pin <= '0'; wait for clk_period*696/2; Pin <= '1'; wait for clk_period*696/2;
Pin <= '0'; wait for clk_period*697/2; Pin <= '1'; wait for clk_period*697/2;
Pin <= '0'; wait for clk_period*698/2; Pin <= '1'; wait for clk_period*698/2;
Pin <= '0'; wait for clk_period*699/2; Pin <= '1'; wait for clk_period*699/2;
Pin <= '0'; wait for clk_period*700/2; Pin <= '1'; wait for clk_period*700/2;
Pin <= '0'; wait for clk_period*701/2; Pin <= '1'; wait for clk_period*701/2;
Pin <= '0'; wait for clk_period*702/2; Pin <= '1'; wait for clk_period*702/2;
Pin <= '0'; wait for clk_period*703/2; Pin <= '1'; wait for clk_period*703/2;
Pin <= '0'; wait for clk_period*704/2; Pin <= '1'; wait for clk_period*704/2;
Pin <= '0'; wait for clk_period*705/2; Pin <= '1'; wait for clk_period*705/2;
Pin <= '0'; wait for clk_period*706/2; Pin <= '1'; wait for clk_period*706/2;
Pin <= '0'; wait for clk_period*707/2; Pin <= '1'; wait for clk_period*707/2;
Pin <= '0'; wait for clk_period*708/2; Pin <= '1'; wait for clk_period*708/2;
Pin <= '0'; wait for clk_period*709/2; Pin <= '1'; wait for clk_period*709/2;
Pin <= '0'; wait for clk_period*710/2; Pin <= '1'; wait for clk_period*710/2;
Pin <= '0'; wait for clk_period*711/2; Pin <= '1'; wait for clk_period*711/2;
Pin <= '0'; wait for clk_period*712/2; Pin <= '1'; wait for clk_period*712/2;
Pin <= '0'; wait for clk_period*713/2; Pin <= '1'; wait for clk_period*713/2;
Pin <= '0'; wait for clk_period*714/2; Pin <= '1'; wait for clk_period*714/2;
Pin <= '0'; wait for clk_period*715/2; Pin <= '1'; wait for clk_period*715/2;
Pin <= '0'; wait for clk_period*716/2; Pin <= '1'; wait for clk_period*716/2;
Pin <= '0'; wait for clk_period*717/2; Pin <= '1'; wait for clk_period*717/2;
Pin <= '0'; wait for clk_period*718/2; Pin <= '1'; wait for clk_period*718/2;
Pin <= '0'; wait for clk_period*719/2; Pin <= '1'; wait for clk_period*719/2;
Pin <= '0'; wait for clk_period*720/2; Pin <= '1'; wait for clk_period*720/2;
Pin <= '0'; wait for clk_period*721/2; Pin <= '1'; wait for clk_period*721/2;
Pin <= '0'; wait for clk_period*722/2; Pin <= '1'; wait for clk_period*722/2;
Pin <= '0'; wait for clk_period*723/2; Pin <= '1'; wait for clk_period*723/2;
Pin <= '0'; wait for clk_period*724/2; Pin <= '1'; wait for clk_period*724/2;
Pin <= '0'; wait for clk_period*725/2; Pin <= '1'; wait for clk_period*725/2;
Pin <= '0'; wait for clk_period*726/2; Pin <= '1'; wait for clk_period*726/2;
Pin <= '0'; wait for clk_period*727/2; Pin <= '1'; wait for clk_period*727/2;
Pin <= '0'; wait for clk_period*728/2; Pin <= '1'; wait for clk_period*728/2;
Pin <= '0'; wait for clk_period*729/2; Pin <= '1'; wait for clk_period*729/2;
Pin <= '0'; wait for clk_period*730/2; Pin <= '1'; wait for clk_period*730/2;
Pin <= '0'; wait for clk_period*731/2; Pin <= '1'; wait for clk_period*731/2;
Pin <= '0'; wait for clk_period*732/2; Pin <= '1'; wait for clk_period*732/2;
Pin <= '0'; wait for clk_period*733/2; Pin <= '1'; wait for clk_period*733/2;
Pin <= '0'; wait for clk_period*734/2; Pin <= '1'; wait for clk_period*734/2;
Pin <= '0'; wait for clk_period*735/2; Pin <= '1'; wait for clk_period*735/2;
Pin <= '0'; wait for clk_period*736/2; Pin <= '1'; wait for clk_period*736/2;
Pin <= '0'; wait for clk_period*737/2; Pin <= '1'; wait for clk_period*737/2;
Pin <= '0'; wait for clk_period*738/2; Pin <= '1'; wait for clk_period*738/2;
Pin <= '0'; wait for clk_period*739/2; Pin <= '1'; wait for clk_period*739/2;
Pin <= '0'; wait for clk_period*740/2; Pin <= '1'; wait for clk_period*740/2;
Pin <= '0'; wait for clk_period*741/2; Pin <= '1'; wait for clk_period*741/2;
Pin <= '0'; wait for clk_period*742/2; Pin <= '1'; wait for clk_period*742/2;
Pin <= '0'; wait for clk_period*743/2; Pin <= '1'; wait for clk_period*743/2;
Pin <= '0'; wait for clk_period*744/2; Pin <= '1'; wait for clk_period*744/2;
Pin <= '0'; wait for clk_period*745/2; Pin <= '1'; wait for clk_period*745/2;
Pin <= '0'; wait for clk_period*746/2; Pin <= '1'; wait for clk_period*746/2;
Pin <= '0'; wait for clk_period*747/2; Pin <= '1'; wait for clk_period*747/2;
Pin <= '0'; wait for clk_period*748/2; Pin <= '1'; wait for clk_period*748/2;
Pin <= '0'; wait for clk_period*749/2; Pin <= '1'; wait for clk_period*749/2;
Pin <= '0'; wait for clk_period*750/2; Pin <= '1'; wait for clk_period*750/2;
Pin <= '0'; wait for clk_period*751/2; Pin <= '1'; wait for clk_period*751/2;
Pin <= '0'; wait for clk_period*752/2; Pin <= '1'; wait for clk_period*752/2;
Pin <= '0'; wait for clk_period*753/2; Pin <= '1'; wait for clk_period*753/2;
Pin <= '0'; wait for clk_period*754/2; Pin <= '1'; wait for clk_period*754/2;
Pin <= '0'; wait for clk_period*755/2; Pin <= '1'; wait for clk_period*755/2;
Pin <= '0'; wait for clk_period*756/2; Pin <= '1'; wait for clk_period*756/2;
Pin <= '0'; wait for clk_period*757/2; Pin <= '1'; wait for clk_period*757/2;
Pin <= '0'; wait for clk_period*758/2; Pin <= '1'; wait for clk_period*758/2;
Pin <= '0'; wait for clk_period*759/2; Pin <= '1'; wait for clk_period*759/2;
Pin <= '0'; wait for clk_period*760/2; Pin <= '1'; wait for clk_period*760/2;
Pin <= '0'; wait for clk_period*761/2; Pin <= '1'; wait for clk_period*761/2;
Pin <= '0'; wait for clk_period*762/2; Pin <= '1'; wait for clk_period*762/2;
Pin <= '0'; wait for clk_period*763/2; Pin <= '1'; wait for clk_period*763/2;
Pin <= '0'; wait for clk_period*764/2; Pin <= '1'; wait for clk_period*764/2;
Pin <= '0'; wait for clk_period*765/2; Pin <= '1'; wait for clk_period*765/2;
Pin <= '0'; wait for clk_period*766/2; Pin <= '1'; wait for clk_period*766/2;
Pin <= '0'; wait for clk_period*767/2; Pin <= '1'; wait for clk_period*767/2;
Pin <= '0'; wait for clk_period*768/2; Pin <= '1'; wait for clk_period*768/2;
Pin <= '0'; wait for clk_period*769/2; Pin <= '1'; wait for clk_period*769/2;
Pin <= '0'; wait for clk_period*770/2; Pin <= '1'; wait for clk_period*770/2;
Pin <= '0'; wait for clk_period*771/2; Pin <= '1'; wait for clk_period*771/2;
Pin <= '0'; wait for clk_period*772/2; Pin <= '1'; wait for clk_period*772/2;
Pin <= '0'; wait for clk_period*773/2; Pin <= '1'; wait for clk_period*773/2;
Pin <= '0'; wait for clk_period*774/2; Pin <= '1'; wait for clk_period*774/2;
Pin <= '0'; wait for clk_period*775/2; Pin <= '1'; wait for clk_period*775/2;
Pin <= '0'; wait for clk_period*776/2; Pin <= '1'; wait for clk_period*776/2;
Pin <= '0'; wait for clk_period*777/2; Pin <= '1'; wait for clk_period*777/2;
Pin <= '0'; wait for clk_period*778/2; Pin <= '1'; wait for clk_period*778/2;
Pin <= '0'; wait for clk_period*779/2; Pin <= '1'; wait for clk_period*779/2;
Pin <= '0'; wait for clk_period*780/2; Pin <= '1'; wait for clk_period*780/2;
Pin <= '0'; wait for clk_period*781/2; Pin <= '1'; wait for clk_period*781/2;
Pin <= '0'; wait for clk_period*782/2; Pin <= '1'; wait for clk_period*782/2;
Pin <= '0'; wait for clk_period*783/2; Pin <= '1'; wait for clk_period*783/2;
Pin <= '0'; wait for clk_period*784/2; Pin <= '1'; wait for clk_period*784/2;
Pin <= '0'; wait for clk_period*785/2; Pin <= '1'; wait for clk_period*785/2;
Pin <= '0'; wait for clk_period*786/2; Pin <= '1'; wait for clk_period*786/2;
Pin <= '0'; wait for clk_period*787/2; Pin <= '1'; wait for clk_period*787/2;
Pin <= '0'; wait for clk_period*788/2; Pin <= '1'; wait for clk_period*788/2;
Pin <= '0'; wait for clk_period*789/2; Pin <= '1'; wait for clk_period*789/2;
Pin <= '0'; wait for clk_period*790/2; Pin <= '1'; wait for clk_period*790/2;
Pin <= '0'; wait for clk_period*791/2; Pin <= '1'; wait for clk_period*791/2;
Pin <= '0'; wait for clk_period*792/2; Pin <= '1'; wait for clk_period*792/2;
Pin <= '0'; wait for clk_period*793/2; Pin <= '1'; wait for clk_period*793/2;
Pin <= '0'; wait for clk_period*794/2; Pin <= '1'; wait for clk_period*794/2;
Pin <= '0'; wait for clk_period*795/2; Pin <= '1'; wait for clk_period*795/2;
Pin <= '0'; wait for clk_period*796/2; Pin <= '1'; wait for clk_period*796/2;
Pin <= '0'; wait for clk_period*797/2; Pin <= '1'; wait for clk_period*797/2;
Pin <= '0'; wait for clk_period*798/2; Pin <= '1'; wait for clk_period*798/2;
Pin <= '0'; wait for clk_period*799/2; Pin <= '1'; wait for clk_period*799/2;
Pin <= '0'; wait for clk_period*800/2; Pin <= '1'; wait for clk_period*800/2;
Pin <= '0'; wait for clk_period*801/2; Pin <= '1'; wait for clk_period*801/2;
Pin <= '0'; wait for clk_period*802/2; Pin <= '1'; wait for clk_period*802/2;
Pin <= '0'; wait for clk_period*803/2; Pin <= '1'; wait for clk_period*803/2;
Pin <= '0'; wait for clk_period*804/2; Pin <= '1'; wait for clk_period*804/2;
Pin <= '0'; wait for clk_period*805/2; Pin <= '1'; wait for clk_period*805/2;
Pin <= '0'; wait for clk_period*806/2; Pin <= '1'; wait for clk_period*806/2;
Pin <= '0'; wait for clk_period*807/2; Pin <= '1'; wait for clk_period*807/2;
Pin <= '0'; wait for clk_period*808/2; Pin <= '1'; wait for clk_period*808/2;
Pin <= '0'; wait for clk_period*809/2; Pin <= '1'; wait for clk_period*809/2;
Pin <= '0'; wait for clk_period*810/2; Pin <= '1'; wait for clk_period*810/2;
Pin <= '0'; wait for clk_period*811/2; Pin <= '1'; wait for clk_period*811/2;
Pin <= '0'; wait for clk_period*812/2; Pin <= '1'; wait for clk_period*812/2;
Pin <= '0'; wait for clk_period*813/2; Pin <= '1'; wait for clk_period*813/2;
Pin <= '0'; wait for clk_period*814/2; Pin <= '1'; wait for clk_period*814/2;
Pin <= '0'; wait for clk_period*815/2; Pin <= '1'; wait for clk_period*815/2;
Pin <= '0'; wait for clk_period*816/2; Pin <= '1'; wait for clk_period*816/2;
Pin <= '0'; wait for clk_period*817/2; Pin <= '1'; wait for clk_period*817/2;
Pin <= '0'; wait for clk_period*818/2; Pin <= '1'; wait for clk_period*818/2;
Pin <= '0'; wait for clk_period*819/2; Pin <= '1'; wait for clk_period*819/2;
Pin <= '0'; wait for clk_period*820/2; Pin <= '1'; wait for clk_period*820/2;
Pin <= '0'; wait for clk_period*821/2; Pin <= '1'; wait for clk_period*821/2;
Pin <= '0'; wait for clk_period*822/2; Pin <= '1'; wait for clk_period*822/2;
Pin <= '0'; wait for clk_period*823/2; Pin <= '1'; wait for clk_period*823/2;
Pin <= '0'; wait for clk_period*824/2; Pin <= '1'; wait for clk_period*824/2;
Pin <= '0'; wait for clk_period*825/2; Pin <= '1'; wait for clk_period*825/2;
Pin <= '0'; wait for clk_period*826/2; Pin <= '1'; wait for clk_period*826/2;
Pin <= '0'; wait for clk_period*827/2; Pin <= '1'; wait for clk_period*827/2;
Pin <= '0'; wait for clk_period*828/2; Pin <= '1'; wait for clk_period*828/2;
Pin <= '0'; wait for clk_period*829/2; Pin <= '1'; wait for clk_period*829/2;
Pin <= '0'; wait for clk_period*830/2; Pin <= '1'; wait for clk_period*830/2;
Pin <= '0'; wait for clk_period*831/2; Pin <= '1'; wait for clk_period*831/2;
Pin <= '0'; wait for clk_period*832/2; Pin <= '1'; wait for clk_period*832/2;
Pin <= '0'; wait for clk_period*833/2; Pin <= '1'; wait for clk_period*833/2;
Pin <= '0'; wait for clk_period*834/2; Pin <= '1'; wait for clk_period*834/2;
Pin <= '0'; wait for clk_period*835/2; Pin <= '1'; wait for clk_period*835/2;
Pin <= '0'; wait for clk_period*836/2; Pin <= '1'; wait for clk_period*836/2;
Pin <= '0'; wait for clk_period*837/2; Pin <= '1'; wait for clk_period*837/2;
Pin <= '0'; wait for clk_period*838/2; Pin <= '1'; wait for clk_period*838/2;
Pin <= '0'; wait for clk_period*839/2; Pin <= '1'; wait for clk_period*839/2;
Pin <= '0'; wait for clk_period*840/2; Pin <= '1'; wait for clk_period*840/2;
Pin <= '0'; wait for clk_period*841/2; Pin <= '1'; wait for clk_period*841/2;
Pin <= '0'; wait for clk_period*842/2; Pin <= '1'; wait for clk_period*842/2;
Pin <= '0'; wait for clk_period*843/2; Pin <= '1'; wait for clk_period*843/2;
Pin <= '0'; wait for clk_period*844/2; Pin <= '1'; wait for clk_period*844/2;
Pin <= '0'; wait for clk_period*845/2; Pin <= '1'; wait for clk_period*845/2;
Pin <= '0'; wait for clk_period*846/2; Pin <= '1'; wait for clk_period*846/2;
Pin <= '0'; wait for clk_period*847/2; Pin <= '1'; wait for clk_period*847/2;
Pin <= '0'; wait for clk_period*848/2; Pin <= '1'; wait for clk_period*848/2;
Pin <= '0'; wait for clk_period*849/2; Pin <= '1'; wait for clk_period*849/2;
Pin <= '0'; wait for clk_period*850/2; Pin <= '1'; wait for clk_period*850/2;
Pin <= '0'; wait for clk_period*851/2; Pin <= '1'; wait for clk_period*851/2;
Pin <= '0'; wait for clk_period*852/2; Pin <= '1'; wait for clk_period*852/2;
Pin <= '0'; wait for clk_period*853/2; Pin <= '1'; wait for clk_period*853/2;
Pin <= '0'; wait for clk_period*854/2; Pin <= '1'; wait for clk_period*854/2;
Pin <= '0'; wait for clk_period*855/2; Pin <= '1'; wait for clk_period*855/2;
Pin <= '0'; wait for clk_period*856/2; Pin <= '1'; wait for clk_period*856/2;
Pin <= '0'; wait for clk_period*857/2; Pin <= '1'; wait for clk_period*857/2;
Pin <= '0'; wait for clk_period*858/2; Pin <= '1'; wait for clk_period*858/2;
Pin <= '0'; wait for clk_period*859/2; Pin <= '1'; wait for clk_period*859/2;
Pin <= '0'; wait for clk_period*860/2; Pin <= '1'; wait for clk_period*860/2;
Pin <= '0'; wait for clk_period*861/2; Pin <= '1'; wait for clk_period*861/2;
Pin <= '0'; wait for clk_period*862/2; Pin <= '1'; wait for clk_period*862/2;
Pin <= '0'; wait for clk_period*863/2; Pin <= '1'; wait for clk_period*863/2;
Pin <= '0'; wait for clk_period*864/2; Pin <= '1'; wait for clk_period*864/2;
Pin <= '0'; wait for clk_period*865/2; Pin <= '1'; wait for clk_period*865/2;
Pin <= '0'; wait for clk_period*866/2; Pin <= '1'; wait for clk_period*866/2;
Pin <= '0'; wait for clk_period*867/2; Pin <= '1'; wait for clk_period*867/2;
Pin <= '0'; wait for clk_period*868/2; Pin <= '1'; wait for clk_period*868/2;
Pin <= '0'; wait for clk_period*869/2; Pin <= '1'; wait for clk_period*869/2;
Pin <= '0'; wait for clk_period*870/2; Pin <= '1'; wait for clk_period*870/2;
Pin <= '0'; wait for clk_period*871/2; Pin <= '1'; wait for clk_period*871/2;
Pin <= '0'; wait for clk_period*872/2; Pin <= '1'; wait for clk_period*872/2;
Pin <= '0'; wait for clk_period*873/2; Pin <= '1'; wait for clk_period*873/2;
Pin <= '0'; wait for clk_period*874/2; Pin <= '1'; wait for clk_period*874/2;
Pin <= '0'; wait for clk_period*875/2; Pin <= '1'; wait for clk_period*875/2;
Pin <= '0'; wait for clk_period*876/2; Pin <= '1'; wait for clk_period*876/2;
Pin <= '0'; wait for clk_period*877/2; Pin <= '1'; wait for clk_period*877/2;
Pin <= '0'; wait for clk_period*878/2; Pin <= '1'; wait for clk_period*878/2;
Pin <= '0'; wait for clk_period*879/2; Pin <= '1'; wait for clk_period*879/2;
Pin <= '0'; wait for clk_period*880/2; Pin <= '1'; wait for clk_period*880/2;
Pin <= '0'; wait for clk_period*881/2; Pin <= '1'; wait for clk_period*881/2;
Pin <= '0'; wait for clk_period*882/2; Pin <= '1'; wait for clk_period*882/2;
Pin <= '0'; wait for clk_period*883/2; Pin <= '1'; wait for clk_period*883/2;
Pin <= '0'; wait for clk_period*884/2; Pin <= '1'; wait for clk_period*884/2;
Pin <= '0'; wait for clk_period*885/2; Pin <= '1'; wait for clk_period*885/2;
Pin <= '0'; wait for clk_period*886/2; Pin <= '1'; wait for clk_period*886/2;
Pin <= '0'; wait for clk_period*887/2; Pin <= '1'; wait for clk_period*887/2;
Pin <= '0'; wait for clk_period*888/2; Pin <= '1'; wait for clk_period*888/2;
Pin <= '0'; wait for clk_period*889/2; Pin <= '1'; wait for clk_period*889/2;
Pin <= '0'; wait for clk_period*890/2; Pin <= '1'; wait for clk_period*890/2;
Pin <= '0'; wait for clk_period*891/2; Pin <= '1'; wait for clk_period*891/2;
Pin <= '0'; wait for clk_period*892/2; Pin <= '1'; wait for clk_period*892/2;
Pin <= '0'; wait for clk_period*893/2; Pin <= '1'; wait for clk_period*893/2;
Pin <= '0'; wait for clk_period*894/2; Pin <= '1'; wait for clk_period*894/2;
Pin <= '0'; wait for clk_period*895/2; Pin <= '1'; wait for clk_period*895/2;
Pin <= '0'; wait for clk_period*896/2; Pin <= '1'; wait for clk_period*896/2;
Pin <= '0'; wait for clk_period*897/2; Pin <= '1'; wait for clk_period*897/2;
Pin <= '0'; wait for clk_period*898/2; Pin <= '1'; wait for clk_period*898/2;
Pin <= '0'; wait for clk_period*899/2; Pin <= '1'; wait for clk_period*899/2;
Pin <= '0'; wait for clk_period*900/2; Pin <= '1'; wait for clk_period*900/2;
Pin <= '0'; wait for clk_period*901/2; Pin <= '1'; wait for clk_period*901/2;
Pin <= '0'; wait for clk_period*902/2; Pin <= '1'; wait for clk_period*902/2;
Pin <= '0'; wait for clk_period*903/2; Pin <= '1'; wait for clk_period*903/2;
Pin <= '0'; wait for clk_period*904/2; Pin <= '1'; wait for clk_period*904/2;
Pin <= '0'; wait for clk_period*905/2; Pin <= '1'; wait for clk_period*905/2;
Pin <= '0'; wait for clk_period*906/2; Pin <= '1'; wait for clk_period*906/2;
Pin <= '0'; wait for clk_period*907/2; Pin <= '1'; wait for clk_period*907/2;
Pin <= '0'; wait for clk_period*908/2; Pin <= '1'; wait for clk_period*908/2;
Pin <= '0'; wait for clk_period*909/2; Pin <= '1'; wait for clk_period*909/2;
Pin <= '0'; wait for clk_period*910/2; Pin <= '1'; wait for clk_period*910/2;
Pin <= '0'; wait for clk_period*911/2; Pin <= '1'; wait for clk_period*911/2;
Pin <= '0'; wait for clk_period*912/2; Pin <= '1'; wait for clk_period*912/2;
Pin <= '0'; wait for clk_period*913/2; Pin <= '1'; wait for clk_period*913/2;
Pin <= '0'; wait for clk_period*914/2; Pin <= '1'; wait for clk_period*914/2;
Pin <= '0'; wait for clk_period*915/2; Pin <= '1'; wait for clk_period*915/2;
Pin <= '0'; wait for clk_period*916/2; Pin <= '1'; wait for clk_period*916/2;
Pin <= '0'; wait for clk_period*917/2; Pin <= '1'; wait for clk_period*917/2;
Pin <= '0'; wait for clk_period*918/2; Pin <= '1'; wait for clk_period*918/2;
Pin <= '0'; wait for clk_period*919/2; Pin <= '1'; wait for clk_period*919/2;
Pin <= '0'; wait for clk_period*920/2; Pin <= '1'; wait for clk_period*920/2;
Pin <= '0'; wait for clk_period*921/2; Pin <= '1'; wait for clk_period*921/2;
Pin <= '0'; wait for clk_period*922/2; Pin <= '1'; wait for clk_period*922/2;
Pin <= '0'; wait for clk_period*923/2; Pin <= '1'; wait for clk_period*923/2;
Pin <= '0'; wait for clk_period*924/2; Pin <= '1'; wait for clk_period*924/2;
Pin <= '0'; wait for clk_period*925/2; Pin <= '1'; wait for clk_period*925/2;
Pin <= '0'; wait for clk_period*926/2; Pin <= '1'; wait for clk_period*926/2;
Pin <= '0'; wait for clk_period*927/2; Pin <= '1'; wait for clk_period*927/2;
Pin <= '0'; wait for clk_period*928/2; Pin <= '1'; wait for clk_period*928/2;
Pin <= '0'; wait for clk_period*929/2; Pin <= '1'; wait for clk_period*929/2;
Pin <= '0'; wait for clk_period*930/2; Pin <= '1'; wait for clk_period*930/2;
Pin <= '0'; wait for clk_period*931/2; Pin <= '1'; wait for clk_period*931/2;
Pin <= '0'; wait for clk_period*932/2; Pin <= '1'; wait for clk_period*932/2;
Pin <= '0'; wait for clk_period*933/2; Pin <= '1'; wait for clk_period*933/2;
Pin <= '0'; wait for clk_period*934/2; Pin <= '1'; wait for clk_period*934/2;
Pin <= '0'; wait for clk_period*935/2; Pin <= '1'; wait for clk_period*935/2;
Pin <= '0'; wait for clk_period*936/2; Pin <= '1'; wait for clk_period*936/2;
Pin <= '0'; wait for clk_period*937/2; Pin <= '1'; wait for clk_period*937/2;
Pin <= '0'; wait for clk_period*938/2; Pin <= '1'; wait for clk_period*938/2;
Pin <= '0'; wait for clk_period*939/2; Pin <= '1'; wait for clk_period*939/2;
Pin <= '0'; wait for clk_period*940/2; Pin <= '1'; wait for clk_period*940/2;
Pin <= '0'; wait for clk_period*941/2; Pin <= '1'; wait for clk_period*941/2;
Pin <= '0'; wait for clk_period*942/2; Pin <= '1'; wait for clk_period*942/2;
Pin <= '0'; wait for clk_period*943/2; Pin <= '1'; wait for clk_period*943/2;
Pin <= '0'; wait for clk_period*944/2; Pin <= '1'; wait for clk_period*944/2;
Pin <= '0'; wait for clk_period*945/2; Pin <= '1'; wait for clk_period*945/2;
Pin <= '0'; wait for clk_period*946/2; Pin <= '1'; wait for clk_period*946/2;
Pin <= '0'; wait for clk_period*947/2; Pin <= '1'; wait for clk_period*947/2;
Pin <= '0'; wait for clk_period*948/2; Pin <= '1'; wait for clk_period*948/2;
Pin <= '0'; wait for clk_period*949/2; Pin <= '1'; wait for clk_period*949/2;
Pin <= '0'; wait for clk_period*950/2; Pin <= '1'; wait for clk_period*950/2;
Pin <= '0'; wait for clk_period*951/2; Pin <= '1'; wait for clk_period*951/2;
Pin <= '0'; wait for clk_period*952/2; Pin <= '1'; wait for clk_period*952/2;
Pin <= '0'; wait for clk_period*953/2; Pin <= '1'; wait for clk_period*953/2;
Pin <= '0'; wait for clk_period*954/2; Pin <= '1'; wait for clk_period*954/2;
Pin <= '0'; wait for clk_period*955/2; Pin <= '1'; wait for clk_period*955/2;
Pin <= '0'; wait for clk_period*956/2; Pin <= '1'; wait for clk_period*956/2;
Pin <= '0'; wait for clk_period*957/2; Pin <= '1'; wait for clk_period*957/2;
Pin <= '0'; wait for clk_period*958/2; Pin <= '1'; wait for clk_period*958/2;
Pin <= '0'; wait for clk_period*959/2; Pin <= '1'; wait for clk_period*959/2;
Pin <= '0'; wait for clk_period*960/2; Pin <= '1'; wait for clk_period*960/2;
Pin <= '0'; wait for clk_period*961/2; Pin <= '1'; wait for clk_period*961/2;
Pin <= '0'; wait for clk_period*962/2; Pin <= '1'; wait for clk_period*962/2;
Pin <= '0'; wait for clk_period*963/2; Pin <= '1'; wait for clk_period*963/2;
Pin <= '0'; wait for clk_period*964/2; Pin <= '1'; wait for clk_period*964/2;
Pin <= '0'; wait for clk_period*965/2; Pin <= '1'; wait for clk_period*965/2;
Pin <= '0'; wait for clk_period*966/2; Pin <= '1'; wait for clk_period*966/2;
Pin <= '0'; wait for clk_period*967/2; Pin <= '1'; wait for clk_period*967/2;
Pin <= '0'; wait for clk_period*968/2; Pin <= '1'; wait for clk_period*968/2;
Pin <= '0'; wait for clk_period*969/2; Pin <= '1'; wait for clk_period*969/2;
Pin <= '0'; wait for clk_period*970/2; Pin <= '1'; wait for clk_period*970/2;
Pin <= '0'; wait for clk_period*971/2; Pin <= '1'; wait for clk_period*971/2;
Pin <= '0'; wait for clk_period*972/2; Pin <= '1'; wait for clk_period*972/2;
Pin <= '0'; wait for clk_period*973/2; Pin <= '1'; wait for clk_period*973/2;
Pin <= '0'; wait for clk_period*974/2; Pin <= '1'; wait for clk_period*974/2;
Pin <= '0'; wait for clk_period*975/2; Pin <= '1'; wait for clk_period*975/2;
Pin <= '0'; wait for clk_period*976/2; Pin <= '1'; wait for clk_period*976/2;
Pin <= '0'; wait for clk_period*977/2; Pin <= '1'; wait for clk_period*977/2;
Pin <= '0'; wait for clk_period*978/2; Pin <= '1'; wait for clk_period*978/2;
Pin <= '0'; wait for clk_period*979/2; Pin <= '1'; wait for clk_period*979/2;
Pin <= '0'; wait for clk_period*980/2; Pin <= '1'; wait for clk_period*980/2;
Pin <= '0'; wait for clk_period*981/2; Pin <= '1'; wait for clk_period*981/2;
Pin <= '0'; wait for clk_period*982/2; Pin <= '1'; wait for clk_period*982/2;
Pin <= '0'; wait for clk_period*983/2; Pin <= '1'; wait for clk_period*983/2;
Pin <= '0'; wait for clk_period*984/2; Pin <= '1'; wait for clk_period*984/2;
Pin <= '0'; wait for clk_period*985/2; Pin <= '1'; wait for clk_period*985/2;
Pin <= '0'; wait for clk_period*986/2; Pin <= '1'; wait for clk_period*986/2;
Pin <= '0'; wait for clk_period*987/2; Pin <= '1'; wait for clk_period*987/2;
Pin <= '0'; wait for clk_period*988/2; Pin <= '1'; wait for clk_period*988/2;
Pin <= '0'; wait for clk_period*989/2; Pin <= '1'; wait for clk_period*989/2;
Pin <= '0'; wait for clk_period*990/2; Pin <= '1'; wait for clk_period*990/2;
Pin <= '0'; wait for clk_period*991/2; Pin <= '1'; wait for clk_period*991/2;
Pin <= '0'; wait for clk_period*992/2; Pin <= '1'; wait for clk_period*992/2;
Pin <= '0'; wait for clk_period*993/2; Pin <= '1'; wait for clk_period*993/2;
Pin <= '0'; wait for clk_period*994/2; Pin <= '1'; wait for clk_period*994/2;
Pin <= '0'; wait for clk_period*995/2; Pin <= '1'; wait for clk_period*995/2;
Pin <= '0'; wait for clk_period*996/2; Pin <= '1'; wait for clk_period*996/2;
Pin <= '0'; wait for clk_period*997/2; Pin <= '1'; wait for clk_period*997/2;
Pin <= '0'; wait for clk_period*998/2; Pin <= '1'; wait for clk_period*998/2;
Pin <= '0'; wait for clk_period*999/2; Pin <= '1'; wait for clk_period*999/2;
Pin <= '0'; wait for clk_period*1000/2; Pin <= '1'; wait for clk_period*1000/2;
Pin <= '0'; wait for clk_period*1001/2; Pin <= '1'; wait for clk_period*1001/2;
Pin <= '0'; wait for clk_period*1002/2; Pin <= '1'; wait for clk_period*1002/2;
Pin <= '0'; wait for clk_period*1003/2; Pin <= '1'; wait for clk_period*1003/2;
Pin <= '0'; wait for clk_period*1004/2; Pin <= '1'; wait for clk_period*1004/2;
Pin <= '0'; wait for clk_period*1005/2; Pin <= '1'; wait for clk_period*1005/2;
Pin <= '0'; wait for clk_period*1006/2; Pin <= '1'; wait for clk_period*1006/2;
Pin <= '0'; wait for clk_period*1007/2; Pin <= '1'; wait for clk_period*1007/2;
Pin <= '0'; wait for clk_period*1008/2; Pin <= '1'; wait for clk_period*1008/2;
Pin <= '0'; wait for clk_period*1009/2; Pin <= '1'; wait for clk_period*1009/2;
Pin <= '0'; wait for clk_period*1010/2; Pin <= '1'; wait for clk_period*1010/2;
Pin <= '0'; wait for clk_period*1011/2; Pin <= '1'; wait for clk_period*1011/2;
Pin <= '0'; wait for clk_period*1012/2; Pin <= '1'; wait for clk_period*1012/2;
Pin <= '0'; wait for clk_period*1013/2; Pin <= '1'; wait for clk_period*1013/2;
Pin <= '0'; wait for clk_period*1014/2; Pin <= '1'; wait for clk_period*1014/2;
Pin <= '0'; wait for clk_period*1015/2; Pin <= '1'; wait for clk_period*1015/2;
Pin <= '0'; wait for clk_period*1016/2; Pin <= '1'; wait for clk_period*1016/2;
Pin <= '0'; wait for clk_period*1017/2; Pin <= '1'; wait for clk_period*1017/2;
Pin <= '0'; wait for clk_period*1018/2; Pin <= '1'; wait for clk_period*1018/2;
Pin <= '0'; wait for clk_period*1019/2; Pin <= '1'; wait for clk_period*1019/2;
Pin <= '0'; wait for clk_period*1020/2; Pin <= '1'; wait for clk_period*1020/2;
Pin <= '0'; wait for clk_period*1021/2; Pin <= '1'; wait for clk_period*1021/2;
Pin <= '0'; wait for clk_period*1022/2; Pin <= '1'; wait for clk_period*1022/2;
Pin <= '0'; wait for clk_period*1023/2; Pin <= '1'; wait for clk_period*1023/2;
Pin <= '0'; wait for clk_period*1024/2; Pin <= '1'; wait for clk_period*1024/2;
Pin <= '0'; wait for clk_period*1025/2; Pin <= '1'; wait for clk_period*1025/2;
Pin <= '0'; wait for clk_period*1026/2; Pin <= '1'; wait for clk_period*1026/2;
Pin <= '0'; wait for clk_period*1027/2; Pin <= '1'; wait for clk_period*1027/2;
Pin <= '0'; wait for clk_period*1028/2; Pin <= '1'; wait for clk_period*1028/2;
Pin <= '0'; wait for clk_period*1029/2; Pin <= '1'; wait for clk_period*1029/2;
Pin <= '0'; wait for clk_period*1030/2; Pin <= '1'; wait for clk_period*1030/2;
Pin <= '0'; wait for clk_period*1031/2; Pin <= '1'; wait for clk_period*1031/2;
Pin <= '0'; wait for clk_period*1032/2; Pin <= '1'; wait for clk_period*1032/2;
Pin <= '0'; wait for clk_period*1033/2; Pin <= '1'; wait for clk_period*1033/2;
Pin <= '0'; wait for clk_period*1034/2; Pin <= '1'; wait for clk_period*1034/2;
Pin <= '0'; wait for clk_period*1035/2; Pin <= '1'; wait for clk_period*1035/2;
Pin <= '0'; wait for clk_period*1036/2; Pin <= '1'; wait for clk_period*1036/2;
Pin <= '0'; wait for clk_period*1037/2; Pin <= '1'; wait for clk_period*1037/2;
Pin <= '0'; wait for clk_period*1038/2; Pin <= '1'; wait for clk_period*1038/2;
Pin <= '0'; wait for clk_period*1039/2; Pin <= '1'; wait for clk_period*1039/2;
Pin <= '0'; wait for clk_period*1040/2; Pin <= '1'; wait for clk_period*1040/2;
Pin <= '0'; wait for clk_period*1041/2; Pin <= '1'; wait for clk_period*1041/2;
Pin <= '0'; wait for clk_period*1042/2; Pin <= '1'; wait for clk_period*1042/2;
Pin <= '0'; wait for clk_period*1043/2; Pin <= '1'; wait for clk_period*1043/2;
Pin <= '0'; wait for clk_period*1044/2; Pin <= '1'; wait for clk_period*1044/2;
Pin <= '0'; wait for clk_period*1045/2; Pin <= '1'; wait for clk_period*1045/2;
Pin <= '0'; wait for clk_period*1046/2; Pin <= '1'; wait for clk_period*1046/2;
Pin <= '0'; wait for clk_period*1047/2; Pin <= '1'; wait for clk_period*1047/2;
Pin <= '0'; wait for clk_period*1048/2; Pin <= '1'; wait for clk_period*1048/2;
Pin <= '0'; wait for clk_period*1049/2; Pin <= '1'; wait for clk_period*1049/2;
Pin <= '0'; wait for clk_period*1050/2; Pin <= '1'; wait for clk_period*1050/2;
Pin <= '0'; wait for clk_period*1051/2; Pin <= '1'; wait for clk_period*1051/2;
Pin <= '0'; wait for clk_period*1052/2; Pin <= '1'; wait for clk_period*1052/2;
Pin <= '0'; wait for clk_period*1053/2; Pin <= '1'; wait for clk_period*1053/2;
Pin <= '0'; wait for clk_period*1054/2; Pin <= '1'; wait for clk_period*1054/2;
Pin <= '0'; wait for clk_period*1055/2; Pin <= '1'; wait for clk_period*1055/2;
Pin <= '0'; wait for clk_period*1056/2; Pin <= '1'; wait for clk_period*1056/2;
Pin <= '0'; wait for clk_period*1057/2; Pin <= '1'; wait for clk_period*1057/2;
Pin <= '0'; wait for clk_period*1058/2; Pin <= '1'; wait for clk_period*1058/2;
Pin <= '0'; wait for clk_period*1059/2; Pin <= '1'; wait for clk_period*1059/2;
Pin <= '0'; wait for clk_period*1060/2; Pin <= '1'; wait for clk_period*1060/2;
Pin <= '0'; wait for clk_period*1061/2; Pin <= '1'; wait for clk_period*1061/2;
Pin <= '0'; wait for clk_period*1062/2; Pin <= '1'; wait for clk_period*1062/2;
Pin <= '0'; wait for clk_period*1063/2; Pin <= '1'; wait for clk_period*1063/2;
Pin <= '0'; wait for clk_period*1064/2; Pin <= '1'; wait for clk_period*1064/2;
Pin <= '0'; wait for clk_period*1065/2; Pin <= '1'; wait for clk_period*1065/2;
Pin <= '0'; wait for clk_period*1066/2; Pin <= '1'; wait for clk_period*1066/2;
Pin <= '0'; wait for clk_period*1067/2; Pin <= '1'; wait for clk_period*1067/2;
Pin <= '0'; wait for clk_period*1068/2; Pin <= '1'; wait for clk_period*1068/2;
Pin <= '0'; wait for clk_period*1069/2; Pin <= '1'; wait for clk_period*1069/2;
Pin <= '0'; wait for clk_period*1070/2; Pin <= '1'; wait for clk_period*1070/2;
Pin <= '0'; wait for clk_period*1071/2; Pin <= '1'; wait for clk_period*1071/2;
Pin <= '0'; wait for clk_period*1072/2; Pin <= '1'; wait for clk_period*1072/2;
Pin <= '0'; wait for clk_period*1073/2; Pin <= '1'; wait for clk_period*1073/2;
Pin <= '0'; wait for clk_period*1074/2; Pin <= '1'; wait for clk_period*1074/2;
Pin <= '0'; wait for clk_period*1075/2; Pin <= '1'; wait for clk_period*1075/2;
Pin <= '0'; wait for clk_period*1076/2; Pin <= '1'; wait for clk_period*1076/2;
Pin <= '0'; wait for clk_period*1077/2; Pin <= '1'; wait for clk_period*1077/2;
Pin <= '0'; wait for clk_period*1078/2; Pin <= '1'; wait for clk_period*1078/2;
Pin <= '0'; wait for clk_period*1079/2; Pin <= '1'; wait for clk_period*1079/2;
Pin <= '0'; wait for clk_period*1080/2; Pin <= '1'; wait for clk_period*1080/2;
Pin <= '0'; wait for clk_period*1081/2; Pin <= '1'; wait for clk_period*1081/2;
Pin <= '0'; wait for clk_period*1082/2; Pin <= '1'; wait for clk_period*1082/2;
Pin <= '0'; wait for clk_period*1083/2; Pin <= '1'; wait for clk_period*1083/2;
Pin <= '0'; wait for clk_period*1084/2; Pin <= '1'; wait for clk_period*1084/2;
Pin <= '0'; wait for clk_period*1085/2; Pin <= '1'; wait for clk_period*1085/2;
Pin <= '0'; wait for clk_period*1086/2; Pin <= '1'; wait for clk_period*1086/2;
Pin <= '0'; wait for clk_period*1087/2; Pin <= '1'; wait for clk_period*1087/2;
Pin <= '0'; wait for clk_period*1088/2; Pin <= '1'; wait for clk_period*1088/2;
Pin <= '0'; wait for clk_period*1089/2; Pin <= '1'; wait for clk_period*1089/2;
Pin <= '0'; wait for clk_period*1090/2; Pin <= '1'; wait for clk_period*1090/2;
Pin <= '0'; wait for clk_period*1091/2; Pin <= '1'; wait for clk_period*1091/2;
Pin <= '0'; wait for clk_period*1092/2; Pin <= '1'; wait for clk_period*1092/2;
Pin <= '0'; wait for clk_period*1093/2; Pin <= '1'; wait for clk_period*1093/2;
Pin <= '0'; wait for clk_period*1094/2; Pin <= '1'; wait for clk_period*1094/2;
Pin <= '0'; wait for clk_period*1095/2; Pin <= '1'; wait for clk_period*1095/2;
Pin <= '0'; wait for clk_period*1096/2; Pin <= '1'; wait for clk_period*1096/2;
Pin <= '0'; wait for clk_period*1097/2; Pin <= '1'; wait for clk_period*1097/2;
Pin <= '0'; wait for clk_period*1098/2; Pin <= '1'; wait for clk_period*1098/2;
Pin <= '0'; wait for clk_period*1099/2; Pin <= '1'; wait for clk_period*1099/2;
Pin <= '0'; wait for clk_period*1100/2; Pin <= '1'; wait for clk_period*1100/2;
Pin <= '0'; wait for clk_period*1101/2; Pin <= '1'; wait for clk_period*1101/2;
Pin <= '0'; wait for clk_period*1102/2; Pin <= '1'; wait for clk_period*1102/2;
Pin <= '0'; wait for clk_period*1103/2; Pin <= '1'; wait for clk_period*1103/2;
Pin <= '0'; wait for clk_period*1104/2; Pin <= '1'; wait for clk_period*1104/2;
Pin <= '0'; wait for clk_period*1105/2; Pin <= '1'; wait for clk_period*1105/2;
Pin <= '0'; wait for clk_period*1106/2; Pin <= '1'; wait for clk_period*1106/2;
Pin <= '0'; wait for clk_period*1107/2; Pin <= '1'; wait for clk_period*1107/2;
Pin <= '0'; wait for clk_period*1108/2; Pin <= '1'; wait for clk_period*1108/2;
Pin <= '0'; wait for clk_period*1109/2; Pin <= '1'; wait for clk_period*1109/2;
Pin <= '0'; wait for clk_period*1110/2; Pin <= '1'; wait for clk_period*1110/2;
Pin <= '0'; wait for clk_period*1111/2; Pin <= '1'; wait for clk_period*1111/2;
Pin <= '0'; wait for clk_period*1112/2; Pin <= '1'; wait for clk_period*1112/2;
Pin <= '0'; wait for clk_period*1113/2; Pin <= '1'; wait for clk_period*1113/2;
Pin <= '0'; wait for clk_period*1114/2; Pin <= '1'; wait for clk_period*1114/2;
Pin <= '0'; wait for clk_period*1115/2; Pin <= '1'; wait for clk_period*1115/2;
Pin <= '0'; wait for clk_period*1116/2; Pin <= '1'; wait for clk_period*1116/2;
Pin <= '0'; wait for clk_period*1117/2; Pin <= '1'; wait for clk_period*1117/2;
Pin <= '0'; wait for clk_period*1118/2; Pin <= '1'; wait for clk_period*1118/2;
Pin <= '0'; wait for clk_period*1119/2; Pin <= '1'; wait for clk_period*1119/2;
Pin <= '0'; wait for clk_period*1120/2; Pin <= '1'; wait for clk_period*1120/2;
Pin <= '0'; wait for clk_period*1121/2; Pin <= '1'; wait for clk_period*1121/2;
Pin <= '0'; wait for clk_period*1122/2; Pin <= '1'; wait for clk_period*1122/2;
Pin <= '0'; wait for clk_period*1123/2; Pin <= '1'; wait for clk_period*1123/2;
Pin <= '0'; wait for clk_period*1124/2; Pin <= '1'; wait for clk_period*1124/2;
Pin <= '0'; wait for clk_period*1125/2; Pin <= '1'; wait for clk_period*1125/2;
Pin <= '0'; wait for clk_period*1126/2; Pin <= '1'; wait for clk_period*1126/2;
Pin <= '0'; wait for clk_period*1127/2; Pin <= '1'; wait for clk_period*1127/2;
Pin <= '0'; wait for clk_period*1128/2; Pin <= '1'; wait for clk_period*1128/2;
Pin <= '0'; wait for clk_period*1129/2; Pin <= '1'; wait for clk_period*1129/2;
Pin <= '0'; wait for clk_period*1130/2; Pin <= '1'; wait for clk_period*1130/2;
Pin <= '0'; wait for clk_period*1131/2; Pin <= '1'; wait for clk_period*1131/2;
Pin <= '0'; wait for clk_period*1132/2; Pin <= '1'; wait for clk_period*1132/2;
Pin <= '0'; wait for clk_period*1133/2; Pin <= '1'; wait for clk_period*1133/2;
Pin <= '0'; wait for clk_period*1134/2; Pin <= '1'; wait for clk_period*1134/2;
Pin <= '0'; wait for clk_period*1135/2; Pin <= '1'; wait for clk_period*1135/2;
Pin <= '0'; wait for clk_period*1136/2; Pin <= '1'; wait for clk_period*1136/2;
Pin <= '0'; wait for clk_period*1137/2; Pin <= '1'; wait for clk_period*1137/2;
Pin <= '0'; wait for clk_period*1138/2; Pin <= '1'; wait for clk_period*1138/2;
Pin <= '0'; wait for clk_period*1139/2; Pin <= '1'; wait for clk_period*1139/2;
Pin <= '0'; wait for clk_period*1140/2; Pin <= '1'; wait for clk_period*1140/2;
Pin <= '0'; wait for clk_period*1141/2; Pin <= '1'; wait for clk_period*1141/2;
Pin <= '0'; wait for clk_period*1142/2; Pin <= '1'; wait for clk_period*1142/2;
Pin <= '0'; wait for clk_period*1143/2; Pin <= '1'; wait for clk_period*1143/2;
Pin <= '0'; wait for clk_period*1144/2; Pin <= '1'; wait for clk_period*1144/2;
Pin <= '0'; wait for clk_period*1145/2; Pin <= '1'; wait for clk_period*1145/2;
Pin <= '0'; wait for clk_period*1146/2; Pin <= '1'; wait for clk_period*1146/2;
Pin <= '0'; wait for clk_period*1147/2; Pin <= '1'; wait for clk_period*1147/2;
Pin <= '0'; wait for clk_period*1148/2; Pin <= '1'; wait for clk_period*1148/2;
Pin <= '0'; wait for clk_period*1149/2; Pin <= '1'; wait for clk_period*1149/2;
Pin <= '0'; wait for clk_period*1150/2; Pin <= '1'; wait for clk_period*1150/2;
Pin <= '0'; wait for clk_period*1151/2; Pin <= '1'; wait for clk_period*1151/2;
Pin <= '0'; wait for clk_period*1152/2; Pin <= '1'; wait for clk_period*1152/2;
Pin <= '0'; wait for clk_period*1153/2; Pin <= '1'; wait for clk_period*1153/2;
Pin <= '0'; wait for clk_period*1154/2; Pin <= '1'; wait for clk_period*1154/2;
Pin <= '0'; wait for clk_period*1155/2; Pin <= '1'; wait for clk_period*1155/2;
Pin <= '0'; wait for clk_period*1156/2; Pin <= '1'; wait for clk_period*1156/2;
Pin <= '0'; wait for clk_period*1157/2; Pin <= '1'; wait for clk_period*1157/2;
Pin <= '0'; wait for clk_period*1158/2; Pin <= '1'; wait for clk_period*1158/2;
Pin <= '0'; wait for clk_period*1159/2; Pin <= '1'; wait for clk_period*1159/2;
Pin <= '0'; wait for clk_period*1160/2; Pin <= '1'; wait for clk_period*1160/2;
Pin <= '0'; wait for clk_period*1161/2; Pin <= '1'; wait for clk_period*1161/2;
Pin <= '0'; wait for clk_period*1162/2; Pin <= '1'; wait for clk_period*1162/2;
Pin <= '0'; wait for clk_period*1163/2; Pin <= '1'; wait for clk_period*1163/2;
Pin <= '0'; wait for clk_period*1164/2; Pin <= '1'; wait for clk_period*1164/2;
Pin <= '0'; wait for clk_period*1165/2; Pin <= '1'; wait for clk_period*1165/2;
Pin <= '0'; wait for clk_period*1166/2; Pin <= '1'; wait for clk_period*1166/2;
Pin <= '0'; wait for clk_period*1167/2; Pin <= '1'; wait for clk_period*1167/2;
Pin <= '0'; wait for clk_period*1168/2; Pin <= '1'; wait for clk_period*1168/2;
Pin <= '0'; wait for clk_period*1169/2; Pin <= '1'; wait for clk_period*1169/2;
Pin <= '0'; wait for clk_period*1170/2; Pin <= '1'; wait for clk_period*1170/2;
Pin <= '0'; wait for clk_period*1171/2; Pin <= '1'; wait for clk_period*1171/2;
Pin <= '0'; wait for clk_period*1172/2; Pin <= '1'; wait for clk_period*1172/2;
Pin <= '0'; wait for clk_period*1173/2; Pin <= '1'; wait for clk_period*1173/2;
Pin <= '0'; wait for clk_period*1174/2; Pin <= '1'; wait for clk_period*1174/2;
Pin <= '0'; wait for clk_period*1175/2; Pin <= '1'; wait for clk_period*1175/2;
Pin <= '0'; wait for clk_period*1176/2; Pin <= '1'; wait for clk_period*1176/2;
Pin <= '0'; wait for clk_period*1177/2; Pin <= '1'; wait for clk_period*1177/2;
Pin <= '0'; wait for clk_period*1178/2; Pin <= '1'; wait for clk_period*1178/2;
Pin <= '0'; wait for clk_period*1179/2; Pin <= '1'; wait for clk_period*1179/2;
Pin <= '0'; wait for clk_period*1180/2; Pin <= '1'; wait for clk_period*1180/2;
Pin <= '0'; wait for clk_period*1181/2; Pin <= '1'; wait for clk_period*1181/2;
Pin <= '0'; wait for clk_period*1182/2; Pin <= '1'; wait for clk_period*1182/2;
Pin <= '0'; wait for clk_period*1183/2; Pin <= '1'; wait for clk_period*1183/2;
Pin <= '0'; wait for clk_period*1184/2; Pin <= '1'; wait for clk_period*1184/2;
Pin <= '0'; wait for clk_period*1185/2; Pin <= '1'; wait for clk_period*1185/2;
Pin <= '0'; wait for clk_period*1186/2; Pin <= '1'; wait for clk_period*1186/2;
Pin <= '0'; wait for clk_period*1187/2; Pin <= '1'; wait for clk_period*1187/2;
Pin <= '0'; wait for clk_period*1188/2; Pin <= '1'; wait for clk_period*1188/2;
Pin <= '0'; wait for clk_period*1189/2; Pin <= '1'; wait for clk_period*1189/2;
Pin <= '0'; wait for clk_period*1190/2; Pin <= '1'; wait for clk_period*1190/2;
Pin <= '0'; wait for clk_period*1191/2; Pin <= '1'; wait for clk_period*1191/2;
Pin <= '0'; wait for clk_period*1192/2; Pin <= '1'; wait for clk_period*1192/2;
Pin <= '0'; wait for clk_period*1193/2; Pin <= '1'; wait for clk_period*1193/2;
Pin <= '0'; wait for clk_period*1194/2; Pin <= '1'; wait for clk_period*1194/2;
Pin <= '0'; wait for clk_period*1195/2; Pin <= '1'; wait for clk_period*1195/2;
Pin <= '0'; wait for clk_period*1196/2; Pin <= '1'; wait for clk_period*1196/2;
Pin <= '0'; wait for clk_period*1197/2; Pin <= '1'; wait for clk_period*1197/2;
Pin <= '0'; wait for clk_period*1198/2; Pin <= '1'; wait for clk_period*1198/2;
Pin <= '0'; wait for clk_period*1199/2; Pin <= '1'; wait for clk_period*1199/2;
Pin <= '0'; wait for clk_period*1200/2; Pin <= '1'; wait for clk_period*1200/2;
Pin <= '0'; wait for clk_period*1201/2; Pin <= '1'; wait for clk_period*1201/2;
Pin <= '0'; wait for clk_period*1202/2; Pin <= '1'; wait for clk_period*1202/2;
Pin <= '0'; wait for clk_period*1203/2; Pin <= '1'; wait for clk_period*1203/2;
Pin <= '0'; wait for clk_period*1204/2; Pin <= '1'; wait for clk_period*1204/2;
Pin <= '0'; wait for clk_period*1205/2; Pin <= '1'; wait for clk_period*1205/2;
Pin <= '0'; wait for clk_period*1206/2; Pin <= '1'; wait for clk_period*1206/2;
Pin <= '0'; wait for clk_period*1207/2; Pin <= '1'; wait for clk_period*1207/2;
Pin <= '0'; wait for clk_period*1208/2; Pin <= '1'; wait for clk_period*1208/2;
Pin <= '0'; wait for clk_period*1209/2; Pin <= '1'; wait for clk_period*1209/2;
Pin <= '0'; wait for clk_period*1210/2; Pin <= '1'; wait for clk_period*1210/2;
Pin <= '0'; wait for clk_period*1211/2; Pin <= '1'; wait for clk_period*1211/2;
Pin <= '0'; wait for clk_period*1212/2; Pin <= '1'; wait for clk_period*1212/2;
Pin <= '0'; wait for clk_period*1213/2; Pin <= '1'; wait for clk_period*1213/2;
Pin <= '0'; wait for clk_period*1214/2; Pin <= '1'; wait for clk_period*1214/2;
Pin <= '0'; wait for clk_period*1215/2; Pin <= '1'; wait for clk_period*1215/2;
Pin <= '0'; wait for clk_period*1216/2; Pin <= '1'; wait for clk_period*1216/2;
Pin <= '0'; wait for clk_period*1217/2; Pin <= '1'; wait for clk_period*1217/2;
Pin <= '0'; wait for clk_period*1218/2; Pin <= '1'; wait for clk_period*1218/2;
Pin <= '0'; wait for clk_period*1219/2; Pin <= '1'; wait for clk_period*1219/2;
Pin <= '0'; wait for clk_period*1220/2; Pin <= '1'; wait for clk_period*1220/2;
Pin <= '0'; wait for clk_period*1221/2; Pin <= '1'; wait for clk_period*1221/2;
Pin <= '0'; wait for clk_period*1222/2; Pin <= '1'; wait for clk_period*1222/2;
Pin <= '0'; wait for clk_period*1223/2; Pin <= '1'; wait for clk_period*1223/2;
Pin <= '0'; wait for clk_period*1224/2; Pin <= '1'; wait for clk_period*1224/2;
Pin <= '0'; wait for clk_period*1225/2; Pin <= '1'; wait for clk_period*1225/2;
Pin <= '0'; wait for clk_period*1226/2; Pin <= '1'; wait for clk_period*1226/2;
Pin <= '0'; wait for clk_period*1227/2; Pin <= '1'; wait for clk_period*1227/2;
Pin <= '0'; wait for clk_period*1228/2; Pin <= '1'; wait for clk_period*1228/2;
Pin <= '0'; wait for clk_period*1229/2; Pin <= '1'; wait for clk_period*1229/2;
Pin <= '0'; wait for clk_period*1230/2; Pin <= '1'; wait for clk_period*1230/2;
Pin <= '0'; wait for clk_period*1231/2; Pin <= '1'; wait for clk_period*1231/2;
Pin <= '0'; wait for clk_period*1232/2; Pin <= '1'; wait for clk_period*1232/2;
Pin <= '0'; wait for clk_period*1233/2; Pin <= '1'; wait for clk_period*1233/2;
Pin <= '0'; wait for clk_period*1234/2; Pin <= '1'; wait for clk_period*1234/2;
Pin <= '0'; wait for clk_period*1235/2; Pin <= '1'; wait for clk_period*1235/2;
Pin <= '0'; wait for clk_period*1236/2; Pin <= '1'; wait for clk_period*1236/2;
Pin <= '0'; wait for clk_period*1237/2; Pin <= '1'; wait for clk_period*1237/2;
Pin <= '0'; wait for clk_period*1238/2; Pin <= '1'; wait for clk_period*1238/2;
Pin <= '0'; wait for clk_period*1239/2; Pin <= '1'; wait for clk_period*1239/2;
Pin <= '0'; wait for clk_period*1240/2; Pin <= '1'; wait for clk_period*1240/2;
Pin <= '0'; wait for clk_period*1241/2; Pin <= '1'; wait for clk_period*1241/2;
Pin <= '0'; wait for clk_period*1242/2; Pin <= '1'; wait for clk_period*1242/2;
Pin <= '0'; wait for clk_period*1243/2; Pin <= '1'; wait for clk_period*1243/2;
Pin <= '0'; wait for clk_period*1244/2; Pin <= '1'; wait for clk_period*1244/2;
Pin <= '0'; wait for clk_period*1245/2; Pin <= '1'; wait for clk_period*1245/2;
Pin <= '0'; wait for clk_period*1246/2; Pin <= '1'; wait for clk_period*1246/2;
Pin <= '0'; wait for clk_period*1247/2; Pin <= '1'; wait for clk_period*1247/2;
Pin <= '0'; wait for clk_period*1248/2; Pin <= '1'; wait for clk_period*1248/2;
Pin <= '0'; wait for clk_period*1249/2; Pin <= '1'; wait for clk_period*1249/2;
Pin <= '0'; wait for clk_period*1250/2; Pin <= '1'; wait for clk_period*1250/2;
Pin <= '0'; wait for clk_period*1251/2; Pin <= '1'; wait for clk_period*1251/2;
Pin <= '0'; wait for clk_period*1252/2; Pin <= '1'; wait for clk_period*1252/2;
Pin <= '0'; wait for clk_period*1253/2; Pin <= '1'; wait for clk_period*1253/2;
Pin <= '0'; wait for clk_period*1254/2; Pin <= '1'; wait for clk_period*1254/2;
Pin <= '0'; wait for clk_period*1255/2; Pin <= '1'; wait for clk_period*1255/2;
Pin <= '0'; wait for clk_period*1256/2; Pin <= '1'; wait for clk_period*1256/2;
Pin <= '0'; wait for clk_period*1257/2; Pin <= '1'; wait for clk_period*1257/2;
Pin <= '0'; wait for clk_period*1258/2; Pin <= '1'; wait for clk_period*1258/2;
Pin <= '0'; wait for clk_period*1259/2; Pin <= '1'; wait for clk_period*1259/2;
Pin <= '0'; wait for clk_period*1260/2; Pin <= '1'; wait for clk_period*1260/2;
Pin <= '0'; wait for clk_period*1261/2; Pin <= '1'; wait for clk_period*1261/2;
Pin <= '0'; wait for clk_period*1262/2; Pin <= '1'; wait for clk_period*1262/2;
Pin <= '0'; wait for clk_period*1263/2; Pin <= '1'; wait for clk_period*1263/2;
Pin <= '0'; wait for clk_period*1264/2; Pin <= '1'; wait for clk_period*1264/2;
Pin <= '0'; wait for clk_period*1265/2; Pin <= '1'; wait for clk_period*1265/2;
Pin <= '0'; wait for clk_period*1266/2; Pin <= '1'; wait for clk_period*1266/2;
Pin <= '0'; wait for clk_period*1267/2; Pin <= '1'; wait for clk_period*1267/2;
Pin <= '0'; wait for clk_period*1268/2; Pin <= '1'; wait for clk_period*1268/2;
Pin <= '0'; wait for clk_period*1269/2; Pin <= '1'; wait for clk_period*1269/2;
Pin <= '0'; wait for clk_period*1270/2; Pin <= '1'; wait for clk_period*1270/2;
Pin <= '0'; wait for clk_period*1271/2; Pin <= '1'; wait for clk_period*1271/2;
Pin <= '0'; wait for clk_period*1272/2; Pin <= '1'; wait for clk_period*1272/2;
Pin <= '0'; wait for clk_period*1273/2; Pin <= '1'; wait for clk_period*1273/2;
Pin <= '0'; wait for clk_period*1274/2; Pin <= '1'; wait for clk_period*1274/2;
Pin <= '0'; wait for clk_period*1275/2; Pin <= '1'; wait for clk_period*1275/2;
Pin <= '0'; wait for clk_period*1276/2; Pin <= '1'; wait for clk_period*1276/2;
Pin <= '0'; wait for clk_period*1277/2; Pin <= '1'; wait for clk_period*1277/2;
Pin <= '0'; wait for clk_period*1278/2; Pin <= '1'; wait for clk_period*1278/2;
Pin <= '0'; wait for clk_period*1279/2; Pin <= '1'; wait for clk_period*1279/2;
Pin <= '0'; wait for clk_period*1280/2; Pin <= '1'; wait for clk_period*1280/2;
Pin <= '0'; wait for clk_period*1281/2; Pin <= '1'; wait for clk_period*1281/2;
Pin <= '0'; wait for clk_period*1282/2; Pin <= '1'; wait for clk_period*1282/2;
Pin <= '0'; wait for clk_period*1283/2; Pin <= '1'; wait for clk_period*1283/2;
Pin <= '0'; wait for clk_period*1284/2; Pin <= '1'; wait for clk_period*1284/2;
Pin <= '0'; wait for clk_period*1285/2; Pin <= '1'; wait for clk_period*1285/2;
Pin <= '0'; wait for clk_period*1286/2; Pin <= '1'; wait for clk_period*1286/2;
Pin <= '0'; wait for clk_period*1287/2; Pin <= '1'; wait for clk_period*1287/2;
Pin <= '0'; wait for clk_period*1288/2; Pin <= '1'; wait for clk_period*1288/2;
Pin <= '0'; wait for clk_period*1289/2; Pin <= '1'; wait for clk_period*1289/2;
Pin <= '0'; wait for clk_period*1290/2; Pin <= '1'; wait for clk_period*1290/2;
Pin <= '0'; wait for clk_period*1291/2; Pin <= '1'; wait for clk_period*1291/2;
Pin <= '0'; wait for clk_period*1292/2; Pin <= '1'; wait for clk_period*1292/2;
Pin <= '0'; wait for clk_period*1293/2; Pin <= '1'; wait for clk_period*1293/2;
Pin <= '0'; wait for clk_period*1294/2; Pin <= '1'; wait for clk_period*1294/2;
Pin <= '0'; wait for clk_period*1295/2; Pin <= '1'; wait for clk_period*1295/2;
Pin <= '0'; wait for clk_period*1296/2; Pin <= '1'; wait for clk_period*1296/2;
Pin <= '0'; wait for clk_period*1297/2; Pin <= '1'; wait for clk_period*1297/2;
Pin <= '0'; wait for clk_period*1298/2; Pin <= '1'; wait for clk_period*1298/2;
Pin <= '0'; wait for clk_period*1299/2; Pin <= '1'; wait for clk_period*1299/2;
Pin <= '0'; wait for clk_period*1300/2; Pin <= '1'; wait for clk_period*1300/2;
Pin <= '0'; wait for clk_period*1301/2; Pin <= '1'; wait for clk_period*1301/2;
Pin <= '0'; wait for clk_period*1302/2; Pin <= '1'; wait for clk_period*1302/2;
Pin <= '0'; wait for clk_period*1303/2; Pin <= '1'; wait for clk_period*1303/2;
Pin <= '0'; wait for clk_period*1304/2; Pin <= '1'; wait for clk_period*1304/2;
Pin <= '0'; wait for clk_period*1305/2; Pin <= '1'; wait for clk_period*1305/2;
Pin <= '0'; wait for clk_period*1306/2; Pin <= '1'; wait for clk_period*1306/2;
Pin <= '0'; wait for clk_period*1307/2; Pin <= '1'; wait for clk_period*1307/2;
Pin <= '0'; wait for clk_period*1308/2; Pin <= '1'; wait for clk_period*1308/2;
Pin <= '0'; wait for clk_period*1309/2; Pin <= '1'; wait for clk_period*1309/2;
Pin <= '0'; wait for clk_period*1310/2; Pin <= '1'; wait for clk_period*1310/2;
Pin <= '0'; wait for clk_period*1311/2; Pin <= '1'; wait for clk_period*1311/2;
Pin <= '0'; wait for clk_period*1312/2; Pin <= '1'; wait for clk_period*1312/2;
Pin <= '0'; wait for clk_period*1313/2; Pin <= '1'; wait for clk_period*1313/2;
Pin <= '0'; wait for clk_period*1314/2; Pin <= '1'; wait for clk_period*1314/2;
Pin <= '0'; wait for clk_period*1315/2; Pin <= '1'; wait for clk_period*1315/2;
Pin <= '0'; wait for clk_period*1316/2; Pin <= '1'; wait for clk_period*1316/2;
Pin <= '0'; wait for clk_period*1317/2; Pin <= '1'; wait for clk_period*1317/2;
Pin <= '0'; wait for clk_period*1318/2; Pin <= '1'; wait for clk_period*1318/2;
Pin <= '0'; wait for clk_period*1319/2; Pin <= '1'; wait for clk_period*1319/2;
Pin <= '0'; wait for clk_period*1320/2; Pin <= '1'; wait for clk_period*1320/2;
Pin <= '0'; wait for clk_period*1321/2; Pin <= '1'; wait for clk_period*1321/2;
Pin <= '0'; wait for clk_period*1322/2; Pin <= '1'; wait for clk_period*1322/2;
Pin <= '0'; wait for clk_period*1323/2; Pin <= '1'; wait for clk_period*1323/2;
Pin <= '0'; wait for clk_period*1324/2; Pin <= '1'; wait for clk_period*1324/2;
Pin <= '0'; wait for clk_period*1325/2; Pin <= '1'; wait for clk_period*1325/2;
Pin <= '0'; wait for clk_period*1326/2; Pin <= '1'; wait for clk_period*1326/2;
Pin <= '0'; wait for clk_period*1327/2; Pin <= '1'; wait for clk_period*1327/2;
Pin <= '0'; wait for clk_period*1328/2; Pin <= '1'; wait for clk_period*1328/2;
Pin <= '0'; wait for clk_period*1329/2; Pin <= '1'; wait for clk_period*1329/2;
Pin <= '0'; wait for clk_period*1330/2; Pin <= '1'; wait for clk_period*1330/2;
Pin <= '0'; wait for clk_period*1331/2; Pin <= '1'; wait for clk_period*1331/2;
Pin <= '0'; wait for clk_period*1332/2; Pin <= '1'; wait for clk_period*1332/2;
Pin <= '0'; wait for clk_period*1333/2; Pin <= '1'; wait for clk_period*1333/2;
Pin <= '0'; wait for clk_period*1334/2; Pin <= '1'; wait for clk_period*1334/2;
Pin <= '0'; wait for clk_period*1335/2; Pin <= '1'; wait for clk_period*1335/2;
Pin <= '0'; wait for clk_period*1336/2; Pin <= '1'; wait for clk_period*1336/2;
Pin <= '0'; wait for clk_period*1337/2; Pin <= '1'; wait for clk_period*1337/2;
Pin <= '0'; wait for clk_period*1338/2; Pin <= '1'; wait for clk_period*1338/2;
Pin <= '0'; wait for clk_period*1339/2; Pin <= '1'; wait for clk_period*1339/2;
Pin <= '0'; wait for clk_period*1340/2; Pin <= '1'; wait for clk_period*1340/2;
Pin <= '0'; wait for clk_period*1341/2; Pin <= '1'; wait for clk_period*1341/2;
Pin <= '0'; wait for clk_period*1342/2; Pin <= '1'; wait for clk_period*1342/2;
Pin <= '0'; wait for clk_period*1343/2; Pin <= '1'; wait for clk_period*1343/2;
Pin <= '0'; wait for clk_period*1344/2; Pin <= '1'; wait for clk_period*1344/2;
Pin <= '0'; wait for clk_period*1345/2; Pin <= '1'; wait for clk_period*1345/2;
Pin <= '0'; wait for clk_period*1346/2; Pin <= '1'; wait for clk_period*1346/2;
Pin <= '0'; wait for clk_period*1347/2; Pin <= '1'; wait for clk_period*1347/2;
Pin <= '0'; wait for clk_period*1348/2; Pin <= '1'; wait for clk_period*1348/2;
Pin <= '0'; wait for clk_period*1349/2; Pin <= '1'; wait for clk_period*1349/2;
Pin <= '0'; wait for clk_period*1350/2; Pin <= '1'; wait for clk_period*1350/2;
Pin <= '0'; wait for clk_period*1351/2; Pin <= '1'; wait for clk_period*1351/2;
Pin <= '0'; wait for clk_period*1352/2; Pin <= '1'; wait for clk_period*1352/2;
Pin <= '0'; wait for clk_period*1353/2; Pin <= '1'; wait for clk_period*1353/2;
Pin <= '0'; wait for clk_period*1354/2; Pin <= '1'; wait for clk_period*1354/2;
Pin <= '0'; wait for clk_period*1355/2; Pin <= '1'; wait for clk_period*1355/2;
Pin <= '0'; wait for clk_period*1356/2; Pin <= '1'; wait for clk_period*1356/2;
Pin <= '0'; wait for clk_period*1357/2; Pin <= '1'; wait for clk_period*1357/2;
Pin <= '0'; wait for clk_period*1358/2; Pin <= '1'; wait for clk_period*1358/2;
Pin <= '0'; wait for clk_period*1359/2; Pin <= '1'; wait for clk_period*1359/2;
Pin <= '0'; wait for clk_period*1360/2; Pin <= '1'; wait for clk_period*1360/2;
Pin <= '0'; wait for clk_period*1361/2; Pin <= '1'; wait for clk_period*1361/2;
Pin <= '0'; wait for clk_period*1362/2; Pin <= '1'; wait for clk_period*1362/2;
Pin <= '0'; wait for clk_period*1363/2; Pin <= '1'; wait for clk_period*1363/2;
Pin <= '0'; wait for clk_period*1364/2; Pin <= '1'; wait for clk_period*1364/2;
Pin <= '0'; wait for clk_period*1365/2; Pin <= '1'; wait for clk_period*1365/2;
Pin <= '0'; wait for clk_period*1366/2; Pin <= '1'; wait for clk_period*1366/2;
Pin <= '0'; wait for clk_period*1367/2; Pin <= '1'; wait for clk_period*1367/2;
Pin <= '0'; wait for clk_period*1368/2; Pin <= '1'; wait for clk_period*1368/2;
Pin <= '0'; wait for clk_period*1369/2; Pin <= '1'; wait for clk_period*1369/2;
Pin <= '0'; wait for clk_period*1370/2; Pin <= '1'; wait for clk_period*1370/2;
Pin <= '0'; wait for clk_period*1371/2; Pin <= '1'; wait for clk_period*1371/2;
Pin <= '0'; wait for clk_period*1372/2; Pin <= '1'; wait for clk_period*1372/2;
Pin <= '0'; wait for clk_period*1373/2; Pin <= '1'; wait for clk_period*1373/2;
Pin <= '0'; wait for clk_period*1374/2; Pin <= '1'; wait for clk_period*1374/2;
Pin <= '0'; wait for clk_period*1375/2; Pin <= '1'; wait for clk_period*1375/2;
Pin <= '0'; wait for clk_period*1376/2; Pin <= '1'; wait for clk_period*1376/2;
Pin <= '0'; wait for clk_period*1377/2; Pin <= '1'; wait for clk_period*1377/2;
Pin <= '0'; wait for clk_period*1378/2; Pin <= '1'; wait for clk_period*1378/2;
Pin <= '0'; wait for clk_period*1379/2; Pin <= '1'; wait for clk_period*1379/2;
Pin <= '0'; wait for clk_period*1380/2; Pin <= '1'; wait for clk_period*1380/2;
Pin <= '0'; wait for clk_period*1381/2; Pin <= '1'; wait for clk_period*1381/2;
Pin <= '0'; wait for clk_period*1382/2; Pin <= '1'; wait for clk_period*1382/2;
Pin <= '0'; wait for clk_period*1383/2; Pin <= '1'; wait for clk_period*1383/2;
Pin <= '0'; wait for clk_period*1384/2; Pin <= '1'; wait for clk_period*1384/2;
Pin <= '0'; wait for clk_period*1385/2; Pin <= '1'; wait for clk_period*1385/2;
Pin <= '0'; wait for clk_period*1386/2; Pin <= '1'; wait for clk_period*1386/2;
Pin <= '0'; wait for clk_period*1387/2; Pin <= '1'; wait for clk_period*1387/2;
Pin <= '0'; wait for clk_period*1388/2; Pin <= '1'; wait for clk_period*1388/2;
Pin <= '0'; wait for clk_period*1389/2; Pin <= '1'; wait for clk_period*1389/2;
Pin <= '0'; wait for clk_period*1390/2; Pin <= '1'; wait for clk_period*1390/2;
Pin <= '0'; wait for clk_period*1391/2; Pin <= '1'; wait for clk_period*1391/2;
Pin <= '0'; wait for clk_period*1392/2; Pin <= '1'; wait for clk_period*1392/2;
Pin <= '0'; wait for clk_period*1393/2; Pin <= '1'; wait for clk_period*1393/2;
Pin <= '0'; wait for clk_period*1394/2; Pin <= '1'; wait for clk_period*1394/2;
Pin <= '0'; wait for clk_period*1395/2; Pin <= '1'; wait for clk_period*1395/2;
Pin <= '0'; wait for clk_period*1396/2; Pin <= '1'; wait for clk_period*1396/2;
Pin <= '0'; wait for clk_period*1397/2; Pin <= '1'; wait for clk_period*1397/2;
Pin <= '0'; wait for clk_period*1398/2; Pin <= '1'; wait for clk_period*1398/2;
Pin <= '0'; wait for clk_period*1399/2; Pin <= '1'; wait for clk_period*1399/2;
Pin <= '0'; wait for clk_period*1400/2; Pin <= '1'; wait for clk_period*1400/2;
Pin <= '0'; wait for clk_period*1401/2; Pin <= '1'; wait for clk_period*1401/2;
Pin <= '0'; wait for clk_period*1402/2; Pin <= '1'; wait for clk_period*1402/2;
Pin <= '0'; wait for clk_period*1403/2; Pin <= '1'; wait for clk_period*1403/2;
Pin <= '0'; wait for clk_period*1404/2; Pin <= '1'; wait for clk_period*1404/2;
Pin <= '0'; wait for clk_period*1405/2; Pin <= '1'; wait for clk_period*1405/2;
Pin <= '0'; wait for clk_period*1406/2; Pin <= '1'; wait for clk_period*1406/2;
Pin <= '0'; wait for clk_period*1407/2; Pin <= '1'; wait for clk_period*1407/2;
Pin <= '0'; wait for clk_period*1408/2; Pin <= '1'; wait for clk_period*1408/2;
Pin <= '0'; wait for clk_period*1409/2; Pin <= '1'; wait for clk_period*1409/2;
Pin <= '0'; wait for clk_period*1410/2; Pin <= '1'; wait for clk_period*1410/2;
Pin <= '0'; wait for clk_period*1411/2; Pin <= '1'; wait for clk_period*1411/2;
Pin <= '0'; wait for clk_period*1412/2; Pin <= '1'; wait for clk_period*1412/2;
Pin <= '0'; wait for clk_period*1413/2; Pin <= '1'; wait for clk_period*1413/2;
Pin <= '0'; wait for clk_period*1414/2; Pin <= '1'; wait for clk_period*1414/2;
Pin <= '0'; wait for clk_period*1415/2; Pin <= '1'; wait for clk_period*1415/2;
Pin <= '0'; wait for clk_period*1416/2; Pin <= '1'; wait for clk_period*1416/2;
Pin <= '0'; wait for clk_period*1417/2; Pin <= '1'; wait for clk_period*1417/2;
Pin <= '0'; wait for clk_period*1418/2; Pin <= '1'; wait for clk_period*1418/2;
Pin <= '0'; wait for clk_period*1419/2; Pin <= '1'; wait for clk_period*1419/2;
Pin <= '0'; wait for clk_period*1420/2; Pin <= '1'; wait for clk_period*1420/2;
Pin <= '0'; wait for clk_period*1421/2; Pin <= '1'; wait for clk_period*1421/2;
Pin <= '0'; wait for clk_period*1422/2; Pin <= '1'; wait for clk_period*1422/2;
Pin <= '0'; wait for clk_period*1423/2; Pin <= '1'; wait for clk_period*1423/2;
Pin <= '0'; wait for clk_period*1424/2; Pin <= '1'; wait for clk_period*1424/2;
Pin <= '0'; wait for clk_period*1425/2; Pin <= '1'; wait for clk_period*1425/2;
Pin <= '0'; wait for clk_period*1426/2; Pin <= '1'; wait for clk_period*1426/2;
Pin <= '0'; wait for clk_period*1427/2; Pin <= '1'; wait for clk_period*1427/2;
Pin <= '0'; wait for clk_period*1428/2; Pin <= '1'; wait for clk_period*1428/2;
Pin <= '0'; wait for clk_period*1429/2; Pin <= '1'; wait for clk_period*1429/2;
Pin <= '0'; wait for clk_period*1430/2; Pin <= '1'; wait for clk_period*1430/2;
Pin <= '0'; wait for clk_period*1431/2; Pin <= '1'; wait for clk_period*1431/2;
Pin <= '0'; wait for clk_period*1432/2; Pin <= '1'; wait for clk_period*1432/2;
Pin <= '0'; wait for clk_period*1433/2; Pin <= '1'; wait for clk_period*1433/2;


   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		delta <= "0000000000000000000000000000000000000000000000000000001000000000";
      wait for clk_period*10;
		rst <= '0';
		wait for clk_period*10;
		rst <= '1';
		wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
