----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 			sergio rivera (srivera (at) ucm.es)
-- 
-- Create Date:    	16:08:08 03/02/2017 
-- Design Name: 
-- Module Name:    	histogram1024 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions:  	
-- Description: 		this HW accepts a binary pulse as input
--							and classifieds it by its time duration
--							in a 1024 bins histogram
--
--							it uses 64bit counters
--
--							the output cable "hist"
--							is the serialized histogram
--
--							the time resolution is T(clk)/2
--							as well as the time base
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments:   this is an initial version
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.ALL;
use IEEE.NUMERIC_STD.ALL;


entity histogram is
    Port ( clk 		: in   STD_LOGIC;
			  rst 		: in   STD_LOGIC;
			  Pin 		: in   STD_LOGIC;
			  delta 		: in   STD_LOGIC_VECTOR ( 63 downto 0 );
			  Pout 		: out  STD_LOGIC;
			  total_time: out  STD_LOGIC_VECTOR ( 63 downto 0 );
           hist 		: out  STD_LOGIC_VECTOR (32767 downto 0)
			 );
end histogram;

architecture Behavioral of histogram is

signal hist0  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist2  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist3  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist4  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist5  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist6  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist7  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist8  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist9  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist10  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist11  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist12  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist13  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist14  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist15  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist16  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist17  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist18  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist19  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist20  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist21  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist22  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist23  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist24  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist25  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist26  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist27  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist28  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist29  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist30  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist31  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist32  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist33  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist34  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist35  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist36  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist37  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist38  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist39  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist40  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist41  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist42  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist43  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist44  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist45  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist46  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist47  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist48  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist49  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist50  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist51  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist52  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist53  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist54  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist55  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist56  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist57  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist58  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist59  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist60  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist61  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist62  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist63  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist64  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist65  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist66  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist67  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist68  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist69  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist70  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist71  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist72  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist73  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist74  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist75  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist76  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist77  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist78  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist79  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist80  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist81  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist82  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist83  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist84  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist85  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist86  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist87  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist88  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist89  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist90  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist91  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist92  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist93  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist94  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist95  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist96  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist97  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist98  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist99  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist100  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist101  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist102  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist103  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist104  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist105  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist106  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist107  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist108  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist109  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist110  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist111  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist112  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist113  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist114  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist115  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist116  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist117  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist118  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist119  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist120  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist121  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist122  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist123  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist124  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist125  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist126  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist127  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist128  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist129  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist130  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist131  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist132  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist133  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist134  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist135  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist136  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist137  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist138  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist139  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist140  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist141  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist142  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist143  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist144  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist145  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist146  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist147  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist148  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist149  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist150  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist151  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist152  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist153  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist154  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist155  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist156  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist157  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist158  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist159  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist160  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist161  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist162  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist163  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist164  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist165  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist166  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist167  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist168  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist169  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist170  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist171  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist172  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist173  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist174  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist175  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist176  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist177  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist178  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist179  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist180  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist181  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist182  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist183  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist184  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist185  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist186  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist187  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist188  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist189  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist190  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist191  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist192  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist193  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist194  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist195  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist196  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist197  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist198  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist199  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist200  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist201  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist202  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist203  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist204  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist205  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist206  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist207  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist208  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist209  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist210  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist211  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist212  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist213  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist214  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist215  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist216  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist217  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist218  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist219  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist220  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist221  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist222  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist223  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist224  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist225  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist226  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist227  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist228  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist229  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist230  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist231  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist232  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist233  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist234  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist235  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist236  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist237  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist238  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist239  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist240  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist241  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist242  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist243  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist244  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist245  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist246  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist247  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist248  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist249  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist250  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist251  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist252  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist253  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist254  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist255  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist256  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist257  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist258  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist259  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist260  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist261  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist262  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist263  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist264  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist265  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist266  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist267  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist268  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist269  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist270  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist271  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist272  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist273  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist274  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist275  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist276  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist277  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist278  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist279  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist280  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist281  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist282  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist283  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist284  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist285  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist286  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist287  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist288  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist289  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist290  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist291  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist292  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist293  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist294  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist295  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist296  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist297  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist298  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist299  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist300  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist301  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist302  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist303  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist304  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist305  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist306  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist307  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist308  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist309  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist310  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist311  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist312  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist313  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist314  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist315  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist316  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist317  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist318  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist319  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist320  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist321  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist322  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist323  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist324  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist325  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist326  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist327  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist328  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist329  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist330  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist331  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist332  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist333  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist334  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist335  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist336  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist337  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist338  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist339  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist340  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist341  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist342  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist343  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist344  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist345  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist346  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist347  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist348  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist349  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist350  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist351  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist352  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist353  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist354  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist355  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist356  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist357  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist358  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist359  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist360  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist361  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist362  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist363  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist364  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist365  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist366  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist367  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist368  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist369  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist370  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist371  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist372  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist373  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist374  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist375  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist376  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist377  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist378  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist379  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist380  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist381  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist382  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist383  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist384  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist385  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist386  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist387  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist388  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist389  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist390  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist391  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist392  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist393  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist394  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist395  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist396  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist397  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist398  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist399  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist400  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist401  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist402  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist403  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist404  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist405  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist406  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist407  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist408  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist409  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist410  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist411  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist412  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist413  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist414  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist415  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist416  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist417  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist418  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist419  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist420  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist421  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist422  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist423  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist424  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist425  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist426  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist427  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist428  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist429  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist430  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist431  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist432  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist433  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist434  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist435  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist436  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist437  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist438  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist439  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist440  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist441  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist442  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist443  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist444  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist445  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist446  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist447  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist448  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist449  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist450  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist451  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist452  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist453  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist454  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist455  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist456  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist457  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist458  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist459  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist460  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist461  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist462  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist463  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist464  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist465  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist466  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist467  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist468  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist469  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist470  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist471  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist472  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist473  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist474  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist475  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist476  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist477  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist478  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist479  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist480  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist481  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist482  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist483  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist484  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist485  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist486  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist487  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist488  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist489  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist490  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist491  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist492  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist493  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist494  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist495  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist496  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist497  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist498  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist499  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist500  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist501  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist502  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist503  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist504  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist505  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist506  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist507  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist508  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist509  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist510  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist511  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist512  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist513  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist514  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist515  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist516  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist517  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist518  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist519  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist520  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist521  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist522  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist523  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist524  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist525  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist526  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist527  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist528  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist529  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist530  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist531  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist532  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist533  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist534  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist535  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist536  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist537  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist538  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist539  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist540  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist541  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist542  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist543  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist544  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist545  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist546  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist547  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist548  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist549  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist550  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist551  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist552  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist553  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist554  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist555  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist556  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist557  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist558  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist559  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist560  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist561  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist562  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist563  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist564  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist565  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist566  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist567  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist568  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist569  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist570  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist571  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist572  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist573  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist574  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist575  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist576  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist577  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist578  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist579  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist580  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist581  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist582  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist583  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist584  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist585  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist586  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist587  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist588  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist589  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist590  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist591  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist592  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist593  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist594  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist595  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist596  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist597  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist598  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist599  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist600  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist601  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist602  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist603  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist604  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist605  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist606  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist607  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist608  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist609  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist610  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist611  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist612  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist613  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist614  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist615  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist616  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist617  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist618  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist619  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist620  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist621  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist622  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist623  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist624  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist625  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist626  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist627  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist628  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist629  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist630  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist631  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist632  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist633  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist634  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist635  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist636  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist637  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist638  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist639  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist640  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist641  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist642  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist643  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist644  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist645  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist646  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist647  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist648  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist649  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist650  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist651  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist652  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist653  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist654  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist655  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist656  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist657  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist658  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist659  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist660  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist661  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist662  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist663  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist664  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist665  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist666  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist667  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist668  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist669  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist670  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist671  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist672  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist673  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist674  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist675  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist676  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist677  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist678  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist679  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist680  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist681  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist682  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist683  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist684  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist685  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist686  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist687  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist688  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist689  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist690  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist691  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist692  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist693  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist694  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist695  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist696  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist697  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist698  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist699  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist700  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist701  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist702  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist703  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist704  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist705  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist706  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist707  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist708  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist709  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist710  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist711  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist712  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist713  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist714  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist715  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist716  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist717  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist718  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist719  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist720  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist721  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist722  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist723  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist724  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist725  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist726  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist727  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist728  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist729  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist730  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist731  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist732  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist733  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist734  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist735  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist736  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist737  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist738  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist739  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist740  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist741  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist742  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist743  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist744  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist745  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist746  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist747  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist748  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist749  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist750  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist751  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist752  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist753  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist754  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist755  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist756  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist757  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist758  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist759  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist760  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist761  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist762  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist763  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist764  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist765  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist766  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist767  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist768  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist769  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist770  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist771  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist772  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist773  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist774  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist775  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist776  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist777  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist778  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist779  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist780  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist781  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist782  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist783  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist784  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist785  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist786  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist787  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist788  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist789  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist790  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist791  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist792  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist793  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist794  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist795  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist796  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist797  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist798  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist799  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist800  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist801  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist802  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist803  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist804  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist805  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist806  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist807  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist808  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist809  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist810  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist811  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist812  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist813  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist814  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist815  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist816  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist817  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist818  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist819  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist820  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist821  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist822  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist823  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist824  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist825  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist826  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist827  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist828  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist829  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist830  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist831  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist832  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist833  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist834  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist835  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist836  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist837  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist838  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist839  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist840  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist841  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist842  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist843  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist844  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist845  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist846  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist847  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist848  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist849  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist850  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist851  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist852  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist853  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist854  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist855  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist856  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist857  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist858  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist859  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist860  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist861  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist862  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist863  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist864  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist865  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist866  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist867  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist868  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist869  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist870  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist871  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist872  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist873  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist874  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist875  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist876  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist877  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist878  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist879  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist880  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist881  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist882  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist883  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist884  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist885  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist886  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist887  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist888  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist889  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist890  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist891  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist892  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist893  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist894  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist895  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist896  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist897  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist898  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist899  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist900  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist901  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist902  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist903  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist904  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist905  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist906  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist907  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist908  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist909  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist910  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist911  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist912  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist913  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist914  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist915  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist916  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist917  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist918  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist919  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist920  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist921  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist922  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist923  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist924  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist925  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist926  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist927  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist928  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist929  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist930  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist931  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist932  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist933  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist934  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist935  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist936  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist937  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist938  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist939  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist940  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist941  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist942  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist943  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist944  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist945  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist946  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist947  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist948  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist949  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist950  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist951  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist952  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist953  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist954  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist955  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist956  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist957  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist958  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist959  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist960  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist961  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist962  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist963  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist964  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist965  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist966  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist967  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist968  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist969  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist970  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist971  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist972  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist973  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist974  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist975  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist976  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist977  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist978  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist979  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist980  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist981  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist982  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist983  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist984  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist985  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist986  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist987  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist988  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist989  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist990  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist991  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist992  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist993  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist994  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist995  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist996  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist997  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist998  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist999  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1000  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1001  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1002  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1003  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1004  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1005  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1006  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1007  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1008  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1009  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1010  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1011  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1012  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1013  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1014  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1015  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1016  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1017  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1018  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1019  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1020  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1021  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1022  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal hist1023  : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal time_gone   : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal time_tmp    : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal time_tmp1   : STD_LOGIC_VECTOR ( 63 downto 0 ) := "0000000000000000000000000000000000000000000000000000000000000000";
signal out_tmp     : STD_LOGIC                        := '0';

begin

process(clk,Pin)
begin
	if rst = '0' then
 		hist0 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist2 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist3 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist4 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist5 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist6 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist7 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist8 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist9 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist10 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist11 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist12 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist13 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist14 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist15 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist16 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist17 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist18 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist19 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist20 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist21 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist22 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist23 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist24 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist25 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist26 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist27 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist28 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist29 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist30 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist31 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist32 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist33 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist34 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist35 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist36 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist37 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist38 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist39 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist40 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist41 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist42 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist43 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist44 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist45 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist46 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist47 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist48 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist49 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist50 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist51 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist52 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist53 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist54 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist55 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist56 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist57 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist58 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist59 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist60 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist61 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist62 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist63 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist64 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist65 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist66 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist67 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist68 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist69 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist70 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist71 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist72 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist73 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist74 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist75 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist76 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist77 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist78 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist79 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist80 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist81 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist82 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist83 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist84 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist85 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist86 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist87 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist88 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist89 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist90 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist91 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist92 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist93 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist94 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist95 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist96 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist97 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist98 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist99 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist100 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist101 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist102 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist103 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist104 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist105 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist106 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist107 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist108 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist109 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist110 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist111 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist112 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist113 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist114 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist115 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist116 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist117 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist118 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist119 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist120 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist121 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist122 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist123 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist124 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist125 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist126 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist127 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist128 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist129 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist130 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist131 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist132 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist133 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist134 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist135 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist136 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist137 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist138 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist139 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist140 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist141 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist142 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist143 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist144 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist145 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist146 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist147 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist148 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist149 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist150 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist151 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist152 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist153 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist154 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist155 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist156 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist157 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist158 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist159 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist160 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist161 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist162 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist163 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist164 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist165 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist166 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist167 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist168 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist169 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist170 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist171 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist172 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist173 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist174 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist175 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist176 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist177 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist178 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist179 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist180 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist181 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist182 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist183 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist184 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist185 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist186 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist187 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist188 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist189 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist190 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist191 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist192 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist193 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist194 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist195 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist196 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist197 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist198 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist199 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist200 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist201 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist202 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist203 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist204 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist205 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist206 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist207 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist208 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist209 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist210 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist211 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist212 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist213 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist214 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist215 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist216 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist217 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist218 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist219 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist220 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist221 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist222 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist223 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist224 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist225 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist226 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist227 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist228 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist229 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist230 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist231 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist232 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist233 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist234 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist235 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist236 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist237 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist238 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist239 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist240 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist241 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist242 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist243 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist244 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist245 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist246 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist247 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist248 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist249 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist250 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist251 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist252 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist253 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist254 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist255 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist256 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist257 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist258 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist259 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist260 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist261 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist262 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist263 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist264 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist265 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist266 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist267 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist268 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist269 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist270 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist271 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist272 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist273 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist274 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist275 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist276 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist277 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist278 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist279 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist280 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist281 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist282 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist283 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist284 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist285 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist286 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist287 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist288 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist289 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist290 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist291 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist292 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist293 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist294 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist295 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist296 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist297 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist298 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist299 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist300 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist301 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist302 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist303 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist304 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist305 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist306 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist307 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist308 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist309 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist310 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist311 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist312 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist313 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist314 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist315 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist316 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist317 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist318 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist319 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist320 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist321 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist322 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist323 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist324 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist325 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist326 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist327 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist328 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist329 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist330 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist331 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist332 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist333 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist334 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist335 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist336 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist337 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist338 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist339 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist340 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist341 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist342 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist343 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist344 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist345 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist346 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist347 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist348 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist349 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist350 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist351 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist352 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist353 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist354 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist355 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist356 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist357 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist358 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist359 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist360 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist361 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist362 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist363 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist364 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist365 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist366 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist367 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist368 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist369 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist370 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist371 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist372 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist373 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist374 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist375 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist376 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist377 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist378 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist379 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist380 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist381 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist382 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist383 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist384 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist385 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist386 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist387 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist388 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist389 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist390 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist391 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist392 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist393 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist394 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist395 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist396 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist397 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist398 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist399 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist400 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist401 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist402 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist403 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist404 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist405 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist406 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist407 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist408 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist409 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist410 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist411 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist412 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist413 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist414 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist415 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist416 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist417 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist418 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist419 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist420 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist421 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist422 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist423 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist424 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist425 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist426 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist427 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist428 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist429 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist430 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist431 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist432 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist433 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist434 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist435 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist436 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist437 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist438 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist439 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist440 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist441 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist442 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist443 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist444 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist445 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist446 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist447 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist448 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist449 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist450 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist451 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist452 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist453 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist454 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist455 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist456 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist457 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist458 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist459 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist460 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist461 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist462 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist463 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist464 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist465 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist466 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist467 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist468 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist469 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist470 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist471 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist472 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist473 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist474 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist475 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist476 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist477 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist478 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist479 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist480 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist481 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist482 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist483 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist484 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist485 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist486 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist487 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist488 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist489 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist490 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist491 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist492 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist493 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist494 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist495 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist496 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist497 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist498 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist499 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist500 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist501 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist502 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist503 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist504 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist505 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist506 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist507 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist508 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist509 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist510 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist511 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist512 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist513 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist514 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist515 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist516 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist517 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist518 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist519 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist520 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist521 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist522 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist523 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist524 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist525 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist526 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist527 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist528 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist529 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist530 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist531 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist532 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist533 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist534 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist535 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist536 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist537 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist538 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist539 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist540 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist541 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist542 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist543 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist544 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist545 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist546 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist547 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist548 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist549 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist550 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist551 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist552 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist553 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist554 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist555 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist556 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist557 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist558 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist559 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist560 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist561 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist562 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist563 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist564 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist565 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist566 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist567 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist568 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist569 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist570 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist571 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist572 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist573 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist574 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist575 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist576 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist577 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist578 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist579 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist580 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist581 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist582 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist583 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist584 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist585 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist586 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist587 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist588 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist589 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist590 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist591 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist592 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist593 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist594 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist595 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist596 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist597 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist598 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist599 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist600 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist601 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist602 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist603 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist604 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist605 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist606 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist607 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist608 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist609 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist610 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist611 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist612 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist613 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist614 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist615 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist616 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist617 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist618 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist619 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist620 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist621 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist622 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist623 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist624 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist625 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist626 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist627 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist628 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist629 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist630 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist631 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist632 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist633 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist634 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist635 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist636 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist637 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist638 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist639 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist640 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist641 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist642 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist643 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist644 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist645 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist646 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist647 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist648 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist649 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist650 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist651 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist652 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist653 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist654 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist655 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist656 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist657 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist658 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist659 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist660 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist661 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist662 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist663 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist664 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist665 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist666 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist667 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist668 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist669 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist670 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist671 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist672 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist673 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist674 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist675 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist676 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist677 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist678 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist679 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist680 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist681 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist682 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist683 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist684 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist685 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist686 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist687 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist688 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist689 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist690 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist691 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist692 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist693 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist694 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist695 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist696 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist697 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist698 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist699 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist700 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist701 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist702 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist703 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist704 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist705 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist706 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist707 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist708 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist709 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist710 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist711 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist712 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist713 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist714 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist715 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist716 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist717 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist718 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist719 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist720 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist721 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist722 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist723 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist724 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist725 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist726 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist727 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist728 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist729 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist730 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist731 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist732 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist733 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist734 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist735 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist736 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist737 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist738 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist739 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist740 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist741 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist742 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist743 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist744 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist745 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist746 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist747 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist748 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist749 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist750 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist751 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist752 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist753 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist754 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist755 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist756 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist757 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist758 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist759 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist760 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist761 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist762 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist763 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist764 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist765 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist766 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist767 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist768 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist769 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist770 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist771 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist772 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist773 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist774 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist775 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist776 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist777 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist778 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist779 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist780 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist781 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist782 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist783 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist784 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist785 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist786 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist787 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist788 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist789 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist790 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist791 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist792 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist793 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist794 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist795 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist796 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist797 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist798 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist799 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist800 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist801 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist802 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist803 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist804 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist805 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist806 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist807 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist808 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist809 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist810 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist811 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist812 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist813 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist814 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist815 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist816 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist817 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist818 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist819 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist820 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist821 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist822 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist823 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist824 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist825 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist826 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist827 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist828 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist829 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist830 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist831 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist832 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist833 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist834 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist835 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist836 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist837 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist838 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist839 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist840 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist841 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist842 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist843 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist844 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist845 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist846 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist847 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist848 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist849 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist850 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist851 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist852 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist853 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist854 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist855 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist856 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist857 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist858 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist859 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist860 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist861 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist862 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist863 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist864 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist865 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist866 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist867 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist868 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist869 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist870 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist871 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist872 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist873 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist874 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist875 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist876 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist877 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist878 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist879 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist880 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist881 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist882 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist883 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist884 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist885 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist886 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist887 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist888 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist889 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist890 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist891 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist892 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist893 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist894 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist895 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist896 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist897 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist898 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist899 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist900 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist901 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist902 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist903 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist904 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist905 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist906 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist907 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist908 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist909 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist910 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist911 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist912 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist913 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist914 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist915 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist916 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist917 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist918 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist919 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist920 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist921 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist922 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist923 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist924 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist925 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist926 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist927 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist928 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist929 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist930 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist931 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist932 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist933 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist934 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist935 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist936 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist937 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist938 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist939 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist940 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist941 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist942 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist943 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist944 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist945 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist946 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist947 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist948 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist949 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist950 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist951 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist952 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist953 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist954 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist955 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist956 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist957 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist958 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist959 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist960 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist961 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist962 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist963 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist964 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist965 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist966 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist967 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist968 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist969 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist970 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist971 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist972 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist973 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist974 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist975 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist976 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist977 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist978 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist979 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist980 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist981 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist982 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist983 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist984 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist985 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist986 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist987 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist988 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist989 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist990 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist991 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist992 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist993 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist994 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist995 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist996 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist997 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist998 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist999 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1000 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1001 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1002 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1003 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1004 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1005 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1006 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1007 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1008 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1009 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1010 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1011 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1012 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1013 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1014 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1015 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1016 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1017 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1018 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1019 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1020 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1021 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1022 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		hist1023 <= "0000000000000000000000000000000000000000000000000000000000000000";
 		time_gone <= "0000000000000000000000000000000000000000000000000000000000000000";
 		time_tmp  <= "0000000000000000000000000000000000000000000000000000000000000000";
 		time_tmp1 <= "0000000000000000000000000000000000000000000000000000000000000000";
		out_tmp   <= '0';
	else
		
	if clk='1' and clk'event then
		time_gone <= time_gone + 1;
	elsif clk='0' and clk'event then
		time_gone <= time_gone + 1;
	end if;
	
	if    Pin'event and time_gone > time_tmp1 and Pin='1' then
		
			time_tmp1 <= time_gone;
				
	elsif Pin'event and time_gone > time_tmp1 and Pin='0' then
	
			out_tmp  <= not out_tmp;
			
			time_tmp <= time_gone-time_tmp1;
		
			if    ((unsigned(time_tmp) > unsigned(delta)*0) and (unsigned(time_tmp) <= unsigned(delta)*1) )  then hist0 <= hist0 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1) and (unsigned(time_tmp) <= unsigned(delta)*2) )  then hist1 <= hist1 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*2) and (unsigned(time_tmp) <= unsigned(delta)*3) )  then hist2 <= hist2 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*3) and (unsigned(time_tmp) <= unsigned(delta)*4) )  then hist3 <= hist3 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*4) and (unsigned(time_tmp) <= unsigned(delta)*5) )  then hist4 <= hist4 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*5) and (unsigned(time_tmp) <= unsigned(delta)*6) )  then hist5 <= hist5 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*6) and (unsigned(time_tmp) <= unsigned(delta)*7) )  then hist6 <= hist6 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*7) and (unsigned(time_tmp) <= unsigned(delta)*8) )  then hist7 <= hist7 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*8) and (unsigned(time_tmp) <= unsigned(delta)*9) )  then hist8 <= hist8 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*9) and (unsigned(time_tmp) <= unsigned(delta)*10) ) then hist9 <= hist9 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*10) and (unsigned(time_tmp) <= unsigned(delta)*11) ) then hist10 <= hist10 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*11) and (unsigned(time_tmp) <= unsigned(delta)*12) ) then hist11 <= hist11 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*12) and (unsigned(time_tmp) <= unsigned(delta)*13) ) then hist12 <= hist12 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*13) and (unsigned(time_tmp) <= unsigned(delta)*14) ) then hist13 <= hist13 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*14) and (unsigned(time_tmp) <= unsigned(delta)*15) ) then hist14 <= hist14 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*15) and (unsigned(time_tmp) <= unsigned(delta)*16) ) then hist15 <= hist15 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*16) and (unsigned(time_tmp) <= unsigned(delta)*17) ) then hist16 <= hist16 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*17) and (unsigned(time_tmp) <= unsigned(delta)*18) ) then hist17 <= hist17 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*18) and (unsigned(time_tmp) <= unsigned(delta)*19) ) then hist18 <= hist18 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*19) and (unsigned(time_tmp) <= unsigned(delta)*20) ) then hist19 <= hist19 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*20) and (unsigned(time_tmp) <= unsigned(delta)*21) ) then hist20 <= hist20 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*21) and (unsigned(time_tmp) <= unsigned(delta)*22) ) then hist21 <= hist21 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*22) and (unsigned(time_tmp) <= unsigned(delta)*23) ) then hist22 <= hist22 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*23) and (unsigned(time_tmp) <= unsigned(delta)*24) ) then hist23 <= hist23 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*24) and (unsigned(time_tmp) <= unsigned(delta)*25) ) then hist24 <= hist24 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*25) and (unsigned(time_tmp) <= unsigned(delta)*26) ) then hist25 <= hist25 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*26) and (unsigned(time_tmp) <= unsigned(delta)*27) ) then hist26 <= hist26 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*27) and (unsigned(time_tmp) <= unsigned(delta)*28) ) then hist27 <= hist27 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*28) and (unsigned(time_tmp) <= unsigned(delta)*29) ) then hist28 <= hist28 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*29) and (unsigned(time_tmp) <= unsigned(delta)*30) ) then hist29 <= hist29 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*30) and (unsigned(time_tmp) <= unsigned(delta)*31) ) then hist30 <= hist30 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*31) and (unsigned(time_tmp) <= unsigned(delta)*32) ) then hist31 <= hist31 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*32) and (unsigned(time_tmp) <= unsigned(delta)*33) ) then hist32 <= hist32 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*33) and (unsigned(time_tmp) <= unsigned(delta)*34) ) then hist33 <= hist33 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*34) and (unsigned(time_tmp) <= unsigned(delta)*35) ) then hist34 <= hist34 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*35) and (unsigned(time_tmp) <= unsigned(delta)*36) ) then hist35 <= hist35 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*36) and (unsigned(time_tmp) <= unsigned(delta)*37) ) then hist36 <= hist36 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*37) and (unsigned(time_tmp) <= unsigned(delta)*38) ) then hist37 <= hist37 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*38) and (unsigned(time_tmp) <= unsigned(delta)*39) ) then hist38 <= hist38 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*39) and (unsigned(time_tmp) <= unsigned(delta)*40) ) then hist39 <= hist39 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*40) and (unsigned(time_tmp) <= unsigned(delta)*41) ) then hist40 <= hist40 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*41) and (unsigned(time_tmp) <= unsigned(delta)*42) ) then hist41 <= hist41 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*42) and (unsigned(time_tmp) <= unsigned(delta)*43) ) then hist42 <= hist42 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*43) and (unsigned(time_tmp) <= unsigned(delta)*44) ) then hist43 <= hist43 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*44) and (unsigned(time_tmp) <= unsigned(delta)*45) ) then hist44 <= hist44 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*45) and (unsigned(time_tmp) <= unsigned(delta)*46) ) then hist45 <= hist45 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*46) and (unsigned(time_tmp) <= unsigned(delta)*47) ) then hist46 <= hist46 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*47) and (unsigned(time_tmp) <= unsigned(delta)*48) ) then hist47 <= hist47 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*48) and (unsigned(time_tmp) <= unsigned(delta)*49) ) then hist48 <= hist48 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*49) and (unsigned(time_tmp) <= unsigned(delta)*50) ) then hist49 <= hist49 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*50) and (unsigned(time_tmp) <= unsigned(delta)*51) ) then hist50 <= hist50 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*51) and (unsigned(time_tmp) <= unsigned(delta)*52) ) then hist51 <= hist51 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*52) and (unsigned(time_tmp) <= unsigned(delta)*53) ) then hist52 <= hist52 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*53) and (unsigned(time_tmp) <= unsigned(delta)*54) ) then hist53 <= hist53 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*54) and (unsigned(time_tmp) <= unsigned(delta)*55) ) then hist54 <= hist54 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*55) and (unsigned(time_tmp) <= unsigned(delta)*56) ) then hist55 <= hist55 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*56) and (unsigned(time_tmp) <= unsigned(delta)*57) ) then hist56 <= hist56 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*57) and (unsigned(time_tmp) <= unsigned(delta)*58) ) then hist57 <= hist57 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*58) and (unsigned(time_tmp) <= unsigned(delta)*59) ) then hist58 <= hist58 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*59) and (unsigned(time_tmp) <= unsigned(delta)*60) ) then hist59 <= hist59 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*60) and (unsigned(time_tmp) <= unsigned(delta)*61) ) then hist60 <= hist60 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*61) and (unsigned(time_tmp) <= unsigned(delta)*62) ) then hist61 <= hist61 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*62) and (unsigned(time_tmp) <= unsigned(delta)*63) ) then hist62 <= hist62 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*63) and (unsigned(time_tmp) <= unsigned(delta)*64) ) then hist63 <= hist63 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*64) and (unsigned(time_tmp) <= unsigned(delta)*65) ) then hist64 <= hist64 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*65) and (unsigned(time_tmp) <= unsigned(delta)*66) ) then hist65 <= hist65 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*66) and (unsigned(time_tmp) <= unsigned(delta)*67) ) then hist66 <= hist66 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*67) and (unsigned(time_tmp) <= unsigned(delta)*68) ) then hist67 <= hist67 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*68) and (unsigned(time_tmp) <= unsigned(delta)*69) ) then hist68 <= hist68 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*69) and (unsigned(time_tmp) <= unsigned(delta)*70) ) then hist69 <= hist69 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*70) and (unsigned(time_tmp) <= unsigned(delta)*71) ) then hist70 <= hist70 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*71) and (unsigned(time_tmp) <= unsigned(delta)*72) ) then hist71 <= hist71 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*72) and (unsigned(time_tmp) <= unsigned(delta)*73) ) then hist72 <= hist72 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*73) and (unsigned(time_tmp) <= unsigned(delta)*74) ) then hist73 <= hist73 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*74) and (unsigned(time_tmp) <= unsigned(delta)*75) ) then hist74 <= hist74 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*75) and (unsigned(time_tmp) <= unsigned(delta)*76) ) then hist75 <= hist75 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*76) and (unsigned(time_tmp) <= unsigned(delta)*77) ) then hist76 <= hist76 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*77) and (unsigned(time_tmp) <= unsigned(delta)*78) ) then hist77 <= hist77 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*78) and (unsigned(time_tmp) <= unsigned(delta)*79) ) then hist78 <= hist78 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*79) and (unsigned(time_tmp) <= unsigned(delta)*80) ) then hist79 <= hist79 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*80) and (unsigned(time_tmp) <= unsigned(delta)*81) ) then hist80 <= hist80 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*81) and (unsigned(time_tmp) <= unsigned(delta)*82) ) then hist81 <= hist81 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*82) and (unsigned(time_tmp) <= unsigned(delta)*83) ) then hist82 <= hist82 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*83) and (unsigned(time_tmp) <= unsigned(delta)*84) ) then hist83 <= hist83 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*84) and (unsigned(time_tmp) <= unsigned(delta)*85) ) then hist84 <= hist84 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*85) and (unsigned(time_tmp) <= unsigned(delta)*86) ) then hist85 <= hist85 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*86) and (unsigned(time_tmp) <= unsigned(delta)*87) ) then hist86 <= hist86 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*87) and (unsigned(time_tmp) <= unsigned(delta)*88) ) then hist87 <= hist87 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*88) and (unsigned(time_tmp) <= unsigned(delta)*89) ) then hist88 <= hist88 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*89) and (unsigned(time_tmp) <= unsigned(delta)*90) ) then hist89 <= hist89 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*90) and (unsigned(time_tmp) <= unsigned(delta)*91) ) then hist90 <= hist90 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*91) and (unsigned(time_tmp) <= unsigned(delta)*92) ) then hist91 <= hist91 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*92) and (unsigned(time_tmp) <= unsigned(delta)*93) ) then hist92 <= hist92 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*93) and (unsigned(time_tmp) <= unsigned(delta)*94) ) then hist93 <= hist93 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*94) and (unsigned(time_tmp) <= unsigned(delta)*95) ) then hist94 <= hist94 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*95) and (unsigned(time_tmp) <= unsigned(delta)*96) ) then hist95 <= hist95 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*96) and (unsigned(time_tmp) <= unsigned(delta)*97) ) then hist96 <= hist96 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*97) and (unsigned(time_tmp) <= unsigned(delta)*98) ) then hist97 <= hist97 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*98) and (unsigned(time_tmp) <= unsigned(delta)*99) ) then hist98 <= hist98 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*99) and (unsigned(time_tmp) <= unsigned(delta)*100) ) then hist99 <= hist99 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*100) and (unsigned(time_tmp) <= unsigned(delta)*101) ) then hist100 <= hist100 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*101) and (unsigned(time_tmp) <= unsigned(delta)*102) ) then hist101 <= hist101 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*102) and (unsigned(time_tmp) <= unsigned(delta)*103) ) then hist102 <= hist102 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*103) and (unsigned(time_tmp) <= unsigned(delta)*104) ) then hist103 <= hist103 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*104) and (unsigned(time_tmp) <= unsigned(delta)*105) ) then hist104 <= hist104 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*105) and (unsigned(time_tmp) <= unsigned(delta)*106) ) then hist105 <= hist105 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*106) and (unsigned(time_tmp) <= unsigned(delta)*107) ) then hist106 <= hist106 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*107) and (unsigned(time_tmp) <= unsigned(delta)*108) ) then hist107 <= hist107 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*108) and (unsigned(time_tmp) <= unsigned(delta)*109) ) then hist108 <= hist108 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*109) and (unsigned(time_tmp) <= unsigned(delta)*110) ) then hist109 <= hist109 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*110) and (unsigned(time_tmp) <= unsigned(delta)*111) ) then hist110 <= hist110 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*111) and (unsigned(time_tmp) <= unsigned(delta)*112) ) then hist111 <= hist111 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*112) and (unsigned(time_tmp) <= unsigned(delta)*113) ) then hist112 <= hist112 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*113) and (unsigned(time_tmp) <= unsigned(delta)*114) ) then hist113 <= hist113 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*114) and (unsigned(time_tmp) <= unsigned(delta)*115) ) then hist114 <= hist114 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*115) and (unsigned(time_tmp) <= unsigned(delta)*116) ) then hist115 <= hist115 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*116) and (unsigned(time_tmp) <= unsigned(delta)*117) ) then hist116 <= hist116 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*117) and (unsigned(time_tmp) <= unsigned(delta)*118) ) then hist117 <= hist117 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*118) and (unsigned(time_tmp) <= unsigned(delta)*119) ) then hist118 <= hist118 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*119) and (unsigned(time_tmp) <= unsigned(delta)*120) ) then hist119 <= hist119 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*120) and (unsigned(time_tmp) <= unsigned(delta)*121) ) then hist120 <= hist120 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*121) and (unsigned(time_tmp) <= unsigned(delta)*122) ) then hist121 <= hist121 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*122) and (unsigned(time_tmp) <= unsigned(delta)*123) ) then hist122 <= hist122 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*123) and (unsigned(time_tmp) <= unsigned(delta)*124) ) then hist123 <= hist123 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*124) and (unsigned(time_tmp) <= unsigned(delta)*125) ) then hist124 <= hist124 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*125) and (unsigned(time_tmp) <= unsigned(delta)*126) ) then hist125 <= hist125 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*126) and (unsigned(time_tmp) <= unsigned(delta)*127) ) then hist126 <= hist126 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*127) and (unsigned(time_tmp) <= unsigned(delta)*128) ) then hist127 <= hist127 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*128) and (unsigned(time_tmp) <= unsigned(delta)*129) ) then hist128 <= hist128 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*129) and (unsigned(time_tmp) <= unsigned(delta)*130) ) then hist129 <= hist129 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*130) and (unsigned(time_tmp) <= unsigned(delta)*131) ) then hist130 <= hist130 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*131) and (unsigned(time_tmp) <= unsigned(delta)*132) ) then hist131 <= hist131 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*132) and (unsigned(time_tmp) <= unsigned(delta)*133) ) then hist132 <= hist132 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*133) and (unsigned(time_tmp) <= unsigned(delta)*134) ) then hist133 <= hist133 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*134) and (unsigned(time_tmp) <= unsigned(delta)*135) ) then hist134 <= hist134 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*135) and (unsigned(time_tmp) <= unsigned(delta)*136) ) then hist135 <= hist135 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*136) and (unsigned(time_tmp) <= unsigned(delta)*137) ) then hist136 <= hist136 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*137) and (unsigned(time_tmp) <= unsigned(delta)*138) ) then hist137 <= hist137 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*138) and (unsigned(time_tmp) <= unsigned(delta)*139) ) then hist138 <= hist138 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*139) and (unsigned(time_tmp) <= unsigned(delta)*140) ) then hist139 <= hist139 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*140) and (unsigned(time_tmp) <= unsigned(delta)*141) ) then hist140 <= hist140 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*141) and (unsigned(time_tmp) <= unsigned(delta)*142) ) then hist141 <= hist141 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*142) and (unsigned(time_tmp) <= unsigned(delta)*143) ) then hist142 <= hist142 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*143) and (unsigned(time_tmp) <= unsigned(delta)*144) ) then hist143 <= hist143 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*144) and (unsigned(time_tmp) <= unsigned(delta)*145) ) then hist144 <= hist144 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*145) and (unsigned(time_tmp) <= unsigned(delta)*146) ) then hist145 <= hist145 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*146) and (unsigned(time_tmp) <= unsigned(delta)*147) ) then hist146 <= hist146 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*147) and (unsigned(time_tmp) <= unsigned(delta)*148) ) then hist147 <= hist147 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*148) and (unsigned(time_tmp) <= unsigned(delta)*149) ) then hist148 <= hist148 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*149) and (unsigned(time_tmp) <= unsigned(delta)*150) ) then hist149 <= hist149 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*150) and (unsigned(time_tmp) <= unsigned(delta)*151) ) then hist150 <= hist150 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*151) and (unsigned(time_tmp) <= unsigned(delta)*152) ) then hist151 <= hist151 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*152) and (unsigned(time_tmp) <= unsigned(delta)*153) ) then hist152 <= hist152 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*153) and (unsigned(time_tmp) <= unsigned(delta)*154) ) then hist153 <= hist153 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*154) and (unsigned(time_tmp) <= unsigned(delta)*155) ) then hist154 <= hist154 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*155) and (unsigned(time_tmp) <= unsigned(delta)*156) ) then hist155 <= hist155 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*156) and (unsigned(time_tmp) <= unsigned(delta)*157) ) then hist156 <= hist156 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*157) and (unsigned(time_tmp) <= unsigned(delta)*158) ) then hist157 <= hist157 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*158) and (unsigned(time_tmp) <= unsigned(delta)*159) ) then hist158 <= hist158 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*159) and (unsigned(time_tmp) <= unsigned(delta)*160) ) then hist159 <= hist159 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*160) and (unsigned(time_tmp) <= unsigned(delta)*161) ) then hist160 <= hist160 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*161) and (unsigned(time_tmp) <= unsigned(delta)*162) ) then hist161 <= hist161 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*162) and (unsigned(time_tmp) <= unsigned(delta)*163) ) then hist162 <= hist162 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*163) and (unsigned(time_tmp) <= unsigned(delta)*164) ) then hist163 <= hist163 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*164) and (unsigned(time_tmp) <= unsigned(delta)*165) ) then hist164 <= hist164 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*165) and (unsigned(time_tmp) <= unsigned(delta)*166) ) then hist165 <= hist165 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*166) and (unsigned(time_tmp) <= unsigned(delta)*167) ) then hist166 <= hist166 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*167) and (unsigned(time_tmp) <= unsigned(delta)*168) ) then hist167 <= hist167 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*168) and (unsigned(time_tmp) <= unsigned(delta)*169) ) then hist168 <= hist168 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*169) and (unsigned(time_tmp) <= unsigned(delta)*170) ) then hist169 <= hist169 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*170) and (unsigned(time_tmp) <= unsigned(delta)*171) ) then hist170 <= hist170 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*171) and (unsigned(time_tmp) <= unsigned(delta)*172) ) then hist171 <= hist171 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*172) and (unsigned(time_tmp) <= unsigned(delta)*173) ) then hist172 <= hist172 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*173) and (unsigned(time_tmp) <= unsigned(delta)*174) ) then hist173 <= hist173 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*174) and (unsigned(time_tmp) <= unsigned(delta)*175) ) then hist174 <= hist174 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*175) and (unsigned(time_tmp) <= unsigned(delta)*176) ) then hist175 <= hist175 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*176) and (unsigned(time_tmp) <= unsigned(delta)*177) ) then hist176 <= hist176 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*177) and (unsigned(time_tmp) <= unsigned(delta)*178) ) then hist177 <= hist177 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*178) and (unsigned(time_tmp) <= unsigned(delta)*179) ) then hist178 <= hist178 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*179) and (unsigned(time_tmp) <= unsigned(delta)*180) ) then hist179 <= hist179 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*180) and (unsigned(time_tmp) <= unsigned(delta)*181) ) then hist180 <= hist180 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*181) and (unsigned(time_tmp) <= unsigned(delta)*182) ) then hist181 <= hist181 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*182) and (unsigned(time_tmp) <= unsigned(delta)*183) ) then hist182 <= hist182 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*183) and (unsigned(time_tmp) <= unsigned(delta)*184) ) then hist183 <= hist183 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*184) and (unsigned(time_tmp) <= unsigned(delta)*185) ) then hist184 <= hist184 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*185) and (unsigned(time_tmp) <= unsigned(delta)*186) ) then hist185 <= hist185 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*186) and (unsigned(time_tmp) <= unsigned(delta)*187) ) then hist186 <= hist186 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*187) and (unsigned(time_tmp) <= unsigned(delta)*188) ) then hist187 <= hist187 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*188) and (unsigned(time_tmp) <= unsigned(delta)*189) ) then hist188 <= hist188 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*189) and (unsigned(time_tmp) <= unsigned(delta)*190) ) then hist189 <= hist189 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*190) and (unsigned(time_tmp) <= unsigned(delta)*191) ) then hist190 <= hist190 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*191) and (unsigned(time_tmp) <= unsigned(delta)*192) ) then hist191 <= hist191 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*192) and (unsigned(time_tmp) <= unsigned(delta)*193) ) then hist192 <= hist192 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*193) and (unsigned(time_tmp) <= unsigned(delta)*194) ) then hist193 <= hist193 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*194) and (unsigned(time_tmp) <= unsigned(delta)*195) ) then hist194 <= hist194 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*195) and (unsigned(time_tmp) <= unsigned(delta)*196) ) then hist195 <= hist195 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*196) and (unsigned(time_tmp) <= unsigned(delta)*197) ) then hist196 <= hist196 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*197) and (unsigned(time_tmp) <= unsigned(delta)*198) ) then hist197 <= hist197 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*198) and (unsigned(time_tmp) <= unsigned(delta)*199) ) then hist198 <= hist198 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*199) and (unsigned(time_tmp) <= unsigned(delta)*200) ) then hist199 <= hist199 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*200) and (unsigned(time_tmp) <= unsigned(delta)*201) ) then hist200 <= hist200 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*201) and (unsigned(time_tmp) <= unsigned(delta)*202) ) then hist201 <= hist201 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*202) and (unsigned(time_tmp) <= unsigned(delta)*203) ) then hist202 <= hist202 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*203) and (unsigned(time_tmp) <= unsigned(delta)*204) ) then hist203 <= hist203 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*204) and (unsigned(time_tmp) <= unsigned(delta)*205) ) then hist204 <= hist204 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*205) and (unsigned(time_tmp) <= unsigned(delta)*206) ) then hist205 <= hist205 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*206) and (unsigned(time_tmp) <= unsigned(delta)*207) ) then hist206 <= hist206 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*207) and (unsigned(time_tmp) <= unsigned(delta)*208) ) then hist207 <= hist207 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*208) and (unsigned(time_tmp) <= unsigned(delta)*209) ) then hist208 <= hist208 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*209) and (unsigned(time_tmp) <= unsigned(delta)*210) ) then hist209 <= hist209 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*210) and (unsigned(time_tmp) <= unsigned(delta)*211) ) then hist210 <= hist210 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*211) and (unsigned(time_tmp) <= unsigned(delta)*212) ) then hist211 <= hist211 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*212) and (unsigned(time_tmp) <= unsigned(delta)*213) ) then hist212 <= hist212 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*213) and (unsigned(time_tmp) <= unsigned(delta)*214) ) then hist213 <= hist213 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*214) and (unsigned(time_tmp) <= unsigned(delta)*215) ) then hist214 <= hist214 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*215) and (unsigned(time_tmp) <= unsigned(delta)*216) ) then hist215 <= hist215 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*216) and (unsigned(time_tmp) <= unsigned(delta)*217) ) then hist216 <= hist216 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*217) and (unsigned(time_tmp) <= unsigned(delta)*218) ) then hist217 <= hist217 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*218) and (unsigned(time_tmp) <= unsigned(delta)*219) ) then hist218 <= hist218 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*219) and (unsigned(time_tmp) <= unsigned(delta)*220) ) then hist219 <= hist219 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*220) and (unsigned(time_tmp) <= unsigned(delta)*221) ) then hist220 <= hist220 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*221) and (unsigned(time_tmp) <= unsigned(delta)*222) ) then hist221 <= hist221 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*222) and (unsigned(time_tmp) <= unsigned(delta)*223) ) then hist222 <= hist222 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*223) and (unsigned(time_tmp) <= unsigned(delta)*224) ) then hist223 <= hist223 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*224) and (unsigned(time_tmp) <= unsigned(delta)*225) ) then hist224 <= hist224 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*225) and (unsigned(time_tmp) <= unsigned(delta)*226) ) then hist225 <= hist225 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*226) and (unsigned(time_tmp) <= unsigned(delta)*227) ) then hist226 <= hist226 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*227) and (unsigned(time_tmp) <= unsigned(delta)*228) ) then hist227 <= hist227 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*228) and (unsigned(time_tmp) <= unsigned(delta)*229) ) then hist228 <= hist228 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*229) and (unsigned(time_tmp) <= unsigned(delta)*230) ) then hist229 <= hist229 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*230) and (unsigned(time_tmp) <= unsigned(delta)*231) ) then hist230 <= hist230 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*231) and (unsigned(time_tmp) <= unsigned(delta)*232) ) then hist231 <= hist231 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*232) and (unsigned(time_tmp) <= unsigned(delta)*233) ) then hist232 <= hist232 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*233) and (unsigned(time_tmp) <= unsigned(delta)*234) ) then hist233 <= hist233 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*234) and (unsigned(time_tmp) <= unsigned(delta)*235) ) then hist234 <= hist234 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*235) and (unsigned(time_tmp) <= unsigned(delta)*236) ) then hist235 <= hist235 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*236) and (unsigned(time_tmp) <= unsigned(delta)*237) ) then hist236 <= hist236 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*237) and (unsigned(time_tmp) <= unsigned(delta)*238) ) then hist237 <= hist237 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*238) and (unsigned(time_tmp) <= unsigned(delta)*239) ) then hist238 <= hist238 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*239) and (unsigned(time_tmp) <= unsigned(delta)*240) ) then hist239 <= hist239 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*240) and (unsigned(time_tmp) <= unsigned(delta)*241) ) then hist240 <= hist240 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*241) and (unsigned(time_tmp) <= unsigned(delta)*242) ) then hist241 <= hist241 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*242) and (unsigned(time_tmp) <= unsigned(delta)*243) ) then hist242 <= hist242 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*243) and (unsigned(time_tmp) <= unsigned(delta)*244) ) then hist243 <= hist243 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*244) and (unsigned(time_tmp) <= unsigned(delta)*245) ) then hist244 <= hist244 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*245) and (unsigned(time_tmp) <= unsigned(delta)*246) ) then hist245 <= hist245 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*246) and (unsigned(time_tmp) <= unsigned(delta)*247) ) then hist246 <= hist246 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*247) and (unsigned(time_tmp) <= unsigned(delta)*248) ) then hist247 <= hist247 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*248) and (unsigned(time_tmp) <= unsigned(delta)*249) ) then hist248 <= hist248 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*249) and (unsigned(time_tmp) <= unsigned(delta)*250) ) then hist249 <= hist249 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*250) and (unsigned(time_tmp) <= unsigned(delta)*251) ) then hist250 <= hist250 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*251) and (unsigned(time_tmp) <= unsigned(delta)*252) ) then hist251 <= hist251 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*252) and (unsigned(time_tmp) <= unsigned(delta)*253) ) then hist252 <= hist252 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*253) and (unsigned(time_tmp) <= unsigned(delta)*254) ) then hist253 <= hist253 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*254) and (unsigned(time_tmp) <= unsigned(delta)*255) ) then hist254 <= hist254 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*255) and (unsigned(time_tmp) <= unsigned(delta)*256) ) then hist255 <= hist255 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*256) and (unsigned(time_tmp) <= unsigned(delta)*257) ) then hist256 <= hist256 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*257) and (unsigned(time_tmp) <= unsigned(delta)*258) ) then hist257 <= hist257 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*258) and (unsigned(time_tmp) <= unsigned(delta)*259) ) then hist258 <= hist258 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*259) and (unsigned(time_tmp) <= unsigned(delta)*260) ) then hist259 <= hist259 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*260) and (unsigned(time_tmp) <= unsigned(delta)*261) ) then hist260 <= hist260 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*261) and (unsigned(time_tmp) <= unsigned(delta)*262) ) then hist261 <= hist261 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*262) and (unsigned(time_tmp) <= unsigned(delta)*263) ) then hist262 <= hist262 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*263) and (unsigned(time_tmp) <= unsigned(delta)*264) ) then hist263 <= hist263 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*264) and (unsigned(time_tmp) <= unsigned(delta)*265) ) then hist264 <= hist264 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*265) and (unsigned(time_tmp) <= unsigned(delta)*266) ) then hist265 <= hist265 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*266) and (unsigned(time_tmp) <= unsigned(delta)*267) ) then hist266 <= hist266 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*267) and (unsigned(time_tmp) <= unsigned(delta)*268) ) then hist267 <= hist267 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*268) and (unsigned(time_tmp) <= unsigned(delta)*269) ) then hist268 <= hist268 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*269) and (unsigned(time_tmp) <= unsigned(delta)*270) ) then hist269 <= hist269 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*270) and (unsigned(time_tmp) <= unsigned(delta)*271) ) then hist270 <= hist270 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*271) and (unsigned(time_tmp) <= unsigned(delta)*272) ) then hist271 <= hist271 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*272) and (unsigned(time_tmp) <= unsigned(delta)*273) ) then hist272 <= hist272 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*273) and (unsigned(time_tmp) <= unsigned(delta)*274) ) then hist273 <= hist273 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*274) and (unsigned(time_tmp) <= unsigned(delta)*275) ) then hist274 <= hist274 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*275) and (unsigned(time_tmp) <= unsigned(delta)*276) ) then hist275 <= hist275 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*276) and (unsigned(time_tmp) <= unsigned(delta)*277) ) then hist276 <= hist276 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*277) and (unsigned(time_tmp) <= unsigned(delta)*278) ) then hist277 <= hist277 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*278) and (unsigned(time_tmp) <= unsigned(delta)*279) ) then hist278 <= hist278 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*279) and (unsigned(time_tmp) <= unsigned(delta)*280) ) then hist279 <= hist279 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*280) and (unsigned(time_tmp) <= unsigned(delta)*281) ) then hist280 <= hist280 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*281) and (unsigned(time_tmp) <= unsigned(delta)*282) ) then hist281 <= hist281 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*282) and (unsigned(time_tmp) <= unsigned(delta)*283) ) then hist282 <= hist282 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*283) and (unsigned(time_tmp) <= unsigned(delta)*284) ) then hist283 <= hist283 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*284) and (unsigned(time_tmp) <= unsigned(delta)*285) ) then hist284 <= hist284 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*285) and (unsigned(time_tmp) <= unsigned(delta)*286) ) then hist285 <= hist285 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*286) and (unsigned(time_tmp) <= unsigned(delta)*287) ) then hist286 <= hist286 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*287) and (unsigned(time_tmp) <= unsigned(delta)*288) ) then hist287 <= hist287 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*288) and (unsigned(time_tmp) <= unsigned(delta)*289) ) then hist288 <= hist288 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*289) and (unsigned(time_tmp) <= unsigned(delta)*290) ) then hist289 <= hist289 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*290) and (unsigned(time_tmp) <= unsigned(delta)*291) ) then hist290 <= hist290 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*291) and (unsigned(time_tmp) <= unsigned(delta)*292) ) then hist291 <= hist291 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*292) and (unsigned(time_tmp) <= unsigned(delta)*293) ) then hist292 <= hist292 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*293) and (unsigned(time_tmp) <= unsigned(delta)*294) ) then hist293 <= hist293 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*294) and (unsigned(time_tmp) <= unsigned(delta)*295) ) then hist294 <= hist294 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*295) and (unsigned(time_tmp) <= unsigned(delta)*296) ) then hist295 <= hist295 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*296) and (unsigned(time_tmp) <= unsigned(delta)*297) ) then hist296 <= hist296 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*297) and (unsigned(time_tmp) <= unsigned(delta)*298) ) then hist297 <= hist297 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*298) and (unsigned(time_tmp) <= unsigned(delta)*299) ) then hist298 <= hist298 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*299) and (unsigned(time_tmp) <= unsigned(delta)*300) ) then hist299 <= hist299 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*300) and (unsigned(time_tmp) <= unsigned(delta)*301) ) then hist300 <= hist300 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*301) and (unsigned(time_tmp) <= unsigned(delta)*302) ) then hist301 <= hist301 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*302) and (unsigned(time_tmp) <= unsigned(delta)*303) ) then hist302 <= hist302 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*303) and (unsigned(time_tmp) <= unsigned(delta)*304) ) then hist303 <= hist303 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*304) and (unsigned(time_tmp) <= unsigned(delta)*305) ) then hist304 <= hist304 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*305) and (unsigned(time_tmp) <= unsigned(delta)*306) ) then hist305 <= hist305 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*306) and (unsigned(time_tmp) <= unsigned(delta)*307) ) then hist306 <= hist306 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*307) and (unsigned(time_tmp) <= unsigned(delta)*308) ) then hist307 <= hist307 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*308) and (unsigned(time_tmp) <= unsigned(delta)*309) ) then hist308 <= hist308 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*309) and (unsigned(time_tmp) <= unsigned(delta)*310) ) then hist309 <= hist309 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*310) and (unsigned(time_tmp) <= unsigned(delta)*311) ) then hist310 <= hist310 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*311) and (unsigned(time_tmp) <= unsigned(delta)*312) ) then hist311 <= hist311 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*312) and (unsigned(time_tmp) <= unsigned(delta)*313) ) then hist312 <= hist312 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*313) and (unsigned(time_tmp) <= unsigned(delta)*314) ) then hist313 <= hist313 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*314) and (unsigned(time_tmp) <= unsigned(delta)*315) ) then hist314 <= hist314 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*315) and (unsigned(time_tmp) <= unsigned(delta)*316) ) then hist315 <= hist315 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*316) and (unsigned(time_tmp) <= unsigned(delta)*317) ) then hist316 <= hist316 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*317) and (unsigned(time_tmp) <= unsigned(delta)*318) ) then hist317 <= hist317 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*318) and (unsigned(time_tmp) <= unsigned(delta)*319) ) then hist318 <= hist318 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*319) and (unsigned(time_tmp) <= unsigned(delta)*320) ) then hist319 <= hist319 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*320) and (unsigned(time_tmp) <= unsigned(delta)*321) ) then hist320 <= hist320 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*321) and (unsigned(time_tmp) <= unsigned(delta)*322) ) then hist321 <= hist321 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*322) and (unsigned(time_tmp) <= unsigned(delta)*323) ) then hist322 <= hist322 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*323) and (unsigned(time_tmp) <= unsigned(delta)*324) ) then hist323 <= hist323 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*324) and (unsigned(time_tmp) <= unsigned(delta)*325) ) then hist324 <= hist324 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*325) and (unsigned(time_tmp) <= unsigned(delta)*326) ) then hist325 <= hist325 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*326) and (unsigned(time_tmp) <= unsigned(delta)*327) ) then hist326 <= hist326 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*327) and (unsigned(time_tmp) <= unsigned(delta)*328) ) then hist327 <= hist327 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*328) and (unsigned(time_tmp) <= unsigned(delta)*329) ) then hist328 <= hist328 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*329) and (unsigned(time_tmp) <= unsigned(delta)*330) ) then hist329 <= hist329 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*330) and (unsigned(time_tmp) <= unsigned(delta)*331) ) then hist330 <= hist330 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*331) and (unsigned(time_tmp) <= unsigned(delta)*332) ) then hist331 <= hist331 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*332) and (unsigned(time_tmp) <= unsigned(delta)*333) ) then hist332 <= hist332 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*333) and (unsigned(time_tmp) <= unsigned(delta)*334) ) then hist333 <= hist333 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*334) and (unsigned(time_tmp) <= unsigned(delta)*335) ) then hist334 <= hist334 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*335) and (unsigned(time_tmp) <= unsigned(delta)*336) ) then hist335 <= hist335 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*336) and (unsigned(time_tmp) <= unsigned(delta)*337) ) then hist336 <= hist336 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*337) and (unsigned(time_tmp) <= unsigned(delta)*338) ) then hist337 <= hist337 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*338) and (unsigned(time_tmp) <= unsigned(delta)*339) ) then hist338 <= hist338 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*339) and (unsigned(time_tmp) <= unsigned(delta)*340) ) then hist339 <= hist339 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*340) and (unsigned(time_tmp) <= unsigned(delta)*341) ) then hist340 <= hist340 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*341) and (unsigned(time_tmp) <= unsigned(delta)*342) ) then hist341 <= hist341 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*342) and (unsigned(time_tmp) <= unsigned(delta)*343) ) then hist342 <= hist342 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*343) and (unsigned(time_tmp) <= unsigned(delta)*344) ) then hist343 <= hist343 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*344) and (unsigned(time_tmp) <= unsigned(delta)*345) ) then hist344 <= hist344 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*345) and (unsigned(time_tmp) <= unsigned(delta)*346) ) then hist345 <= hist345 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*346) and (unsigned(time_tmp) <= unsigned(delta)*347) ) then hist346 <= hist346 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*347) and (unsigned(time_tmp) <= unsigned(delta)*348) ) then hist347 <= hist347 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*348) and (unsigned(time_tmp) <= unsigned(delta)*349) ) then hist348 <= hist348 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*349) and (unsigned(time_tmp) <= unsigned(delta)*350) ) then hist349 <= hist349 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*350) and (unsigned(time_tmp) <= unsigned(delta)*351) ) then hist350 <= hist350 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*351) and (unsigned(time_tmp) <= unsigned(delta)*352) ) then hist351 <= hist351 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*352) and (unsigned(time_tmp) <= unsigned(delta)*353) ) then hist352 <= hist352 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*353) and (unsigned(time_tmp) <= unsigned(delta)*354) ) then hist353 <= hist353 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*354) and (unsigned(time_tmp) <= unsigned(delta)*355) ) then hist354 <= hist354 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*355) and (unsigned(time_tmp) <= unsigned(delta)*356) ) then hist355 <= hist355 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*356) and (unsigned(time_tmp) <= unsigned(delta)*357) ) then hist356 <= hist356 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*357) and (unsigned(time_tmp) <= unsigned(delta)*358) ) then hist357 <= hist357 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*358) and (unsigned(time_tmp) <= unsigned(delta)*359) ) then hist358 <= hist358 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*359) and (unsigned(time_tmp) <= unsigned(delta)*360) ) then hist359 <= hist359 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*360) and (unsigned(time_tmp) <= unsigned(delta)*361) ) then hist360 <= hist360 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*361) and (unsigned(time_tmp) <= unsigned(delta)*362) ) then hist361 <= hist361 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*362) and (unsigned(time_tmp) <= unsigned(delta)*363) ) then hist362 <= hist362 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*363) and (unsigned(time_tmp) <= unsigned(delta)*364) ) then hist363 <= hist363 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*364) and (unsigned(time_tmp) <= unsigned(delta)*365) ) then hist364 <= hist364 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*365) and (unsigned(time_tmp) <= unsigned(delta)*366) ) then hist365 <= hist365 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*366) and (unsigned(time_tmp) <= unsigned(delta)*367) ) then hist366 <= hist366 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*367) and (unsigned(time_tmp) <= unsigned(delta)*368) ) then hist367 <= hist367 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*368) and (unsigned(time_tmp) <= unsigned(delta)*369) ) then hist368 <= hist368 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*369) and (unsigned(time_tmp) <= unsigned(delta)*370) ) then hist369 <= hist369 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*370) and (unsigned(time_tmp) <= unsigned(delta)*371) ) then hist370 <= hist370 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*371) and (unsigned(time_tmp) <= unsigned(delta)*372) ) then hist371 <= hist371 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*372) and (unsigned(time_tmp) <= unsigned(delta)*373) ) then hist372 <= hist372 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*373) and (unsigned(time_tmp) <= unsigned(delta)*374) ) then hist373 <= hist373 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*374) and (unsigned(time_tmp) <= unsigned(delta)*375) ) then hist374 <= hist374 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*375) and (unsigned(time_tmp) <= unsigned(delta)*376) ) then hist375 <= hist375 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*376) and (unsigned(time_tmp) <= unsigned(delta)*377) ) then hist376 <= hist376 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*377) and (unsigned(time_tmp) <= unsigned(delta)*378) ) then hist377 <= hist377 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*378) and (unsigned(time_tmp) <= unsigned(delta)*379) ) then hist378 <= hist378 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*379) and (unsigned(time_tmp) <= unsigned(delta)*380) ) then hist379 <= hist379 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*380) and (unsigned(time_tmp) <= unsigned(delta)*381) ) then hist380 <= hist380 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*381) and (unsigned(time_tmp) <= unsigned(delta)*382) ) then hist381 <= hist381 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*382) and (unsigned(time_tmp) <= unsigned(delta)*383) ) then hist382 <= hist382 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*383) and (unsigned(time_tmp) <= unsigned(delta)*384) ) then hist383 <= hist383 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*384) and (unsigned(time_tmp) <= unsigned(delta)*385) ) then hist384 <= hist384 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*385) and (unsigned(time_tmp) <= unsigned(delta)*386) ) then hist385 <= hist385 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*386) and (unsigned(time_tmp) <= unsigned(delta)*387) ) then hist386 <= hist386 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*387) and (unsigned(time_tmp) <= unsigned(delta)*388) ) then hist387 <= hist387 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*388) and (unsigned(time_tmp) <= unsigned(delta)*389) ) then hist388 <= hist388 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*389) and (unsigned(time_tmp) <= unsigned(delta)*390) ) then hist389 <= hist389 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*390) and (unsigned(time_tmp) <= unsigned(delta)*391) ) then hist390 <= hist390 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*391) and (unsigned(time_tmp) <= unsigned(delta)*392) ) then hist391 <= hist391 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*392) and (unsigned(time_tmp) <= unsigned(delta)*393) ) then hist392 <= hist392 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*393) and (unsigned(time_tmp) <= unsigned(delta)*394) ) then hist393 <= hist393 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*394) and (unsigned(time_tmp) <= unsigned(delta)*395) ) then hist394 <= hist394 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*395) and (unsigned(time_tmp) <= unsigned(delta)*396) ) then hist395 <= hist395 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*396) and (unsigned(time_tmp) <= unsigned(delta)*397) ) then hist396 <= hist396 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*397) and (unsigned(time_tmp) <= unsigned(delta)*398) ) then hist397 <= hist397 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*398) and (unsigned(time_tmp) <= unsigned(delta)*399) ) then hist398 <= hist398 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*399) and (unsigned(time_tmp) <= unsigned(delta)*400) ) then hist399 <= hist399 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*400) and (unsigned(time_tmp) <= unsigned(delta)*401) ) then hist400 <= hist400 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*401) and (unsigned(time_tmp) <= unsigned(delta)*402) ) then hist401 <= hist401 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*402) and (unsigned(time_tmp) <= unsigned(delta)*403) ) then hist402 <= hist402 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*403) and (unsigned(time_tmp) <= unsigned(delta)*404) ) then hist403 <= hist403 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*404) and (unsigned(time_tmp) <= unsigned(delta)*405) ) then hist404 <= hist404 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*405) and (unsigned(time_tmp) <= unsigned(delta)*406) ) then hist405 <= hist405 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*406) and (unsigned(time_tmp) <= unsigned(delta)*407) ) then hist406 <= hist406 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*407) and (unsigned(time_tmp) <= unsigned(delta)*408) ) then hist407 <= hist407 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*408) and (unsigned(time_tmp) <= unsigned(delta)*409) ) then hist408 <= hist408 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*409) and (unsigned(time_tmp) <= unsigned(delta)*410) ) then hist409 <= hist409 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*410) and (unsigned(time_tmp) <= unsigned(delta)*411) ) then hist410 <= hist410 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*411) and (unsigned(time_tmp) <= unsigned(delta)*412) ) then hist411 <= hist411 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*412) and (unsigned(time_tmp) <= unsigned(delta)*413) ) then hist412 <= hist412 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*413) and (unsigned(time_tmp) <= unsigned(delta)*414) ) then hist413 <= hist413 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*414) and (unsigned(time_tmp) <= unsigned(delta)*415) ) then hist414 <= hist414 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*415) and (unsigned(time_tmp) <= unsigned(delta)*416) ) then hist415 <= hist415 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*416) and (unsigned(time_tmp) <= unsigned(delta)*417) ) then hist416 <= hist416 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*417) and (unsigned(time_tmp) <= unsigned(delta)*418) ) then hist417 <= hist417 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*418) and (unsigned(time_tmp) <= unsigned(delta)*419) ) then hist418 <= hist418 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*419) and (unsigned(time_tmp) <= unsigned(delta)*420) ) then hist419 <= hist419 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*420) and (unsigned(time_tmp) <= unsigned(delta)*421) ) then hist420 <= hist420 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*421) and (unsigned(time_tmp) <= unsigned(delta)*422) ) then hist421 <= hist421 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*422) and (unsigned(time_tmp) <= unsigned(delta)*423) ) then hist422 <= hist422 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*423) and (unsigned(time_tmp) <= unsigned(delta)*424) ) then hist423 <= hist423 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*424) and (unsigned(time_tmp) <= unsigned(delta)*425) ) then hist424 <= hist424 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*425) and (unsigned(time_tmp) <= unsigned(delta)*426) ) then hist425 <= hist425 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*426) and (unsigned(time_tmp) <= unsigned(delta)*427) ) then hist426 <= hist426 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*427) and (unsigned(time_tmp) <= unsigned(delta)*428) ) then hist427 <= hist427 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*428) and (unsigned(time_tmp) <= unsigned(delta)*429) ) then hist428 <= hist428 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*429) and (unsigned(time_tmp) <= unsigned(delta)*430) ) then hist429 <= hist429 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*430) and (unsigned(time_tmp) <= unsigned(delta)*431) ) then hist430 <= hist430 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*431) and (unsigned(time_tmp) <= unsigned(delta)*432) ) then hist431 <= hist431 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*432) and (unsigned(time_tmp) <= unsigned(delta)*433) ) then hist432 <= hist432 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*433) and (unsigned(time_tmp) <= unsigned(delta)*434) ) then hist433 <= hist433 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*434) and (unsigned(time_tmp) <= unsigned(delta)*435) ) then hist434 <= hist434 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*435) and (unsigned(time_tmp) <= unsigned(delta)*436) ) then hist435 <= hist435 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*436) and (unsigned(time_tmp) <= unsigned(delta)*437) ) then hist436 <= hist436 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*437) and (unsigned(time_tmp) <= unsigned(delta)*438) ) then hist437 <= hist437 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*438) and (unsigned(time_tmp) <= unsigned(delta)*439) ) then hist438 <= hist438 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*439) and (unsigned(time_tmp) <= unsigned(delta)*440) ) then hist439 <= hist439 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*440) and (unsigned(time_tmp) <= unsigned(delta)*441) ) then hist440 <= hist440 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*441) and (unsigned(time_tmp) <= unsigned(delta)*442) ) then hist441 <= hist441 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*442) and (unsigned(time_tmp) <= unsigned(delta)*443) ) then hist442 <= hist442 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*443) and (unsigned(time_tmp) <= unsigned(delta)*444) ) then hist443 <= hist443 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*444) and (unsigned(time_tmp) <= unsigned(delta)*445) ) then hist444 <= hist444 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*445) and (unsigned(time_tmp) <= unsigned(delta)*446) ) then hist445 <= hist445 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*446) and (unsigned(time_tmp) <= unsigned(delta)*447) ) then hist446 <= hist446 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*447) and (unsigned(time_tmp) <= unsigned(delta)*448) ) then hist447 <= hist447 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*448) and (unsigned(time_tmp) <= unsigned(delta)*449) ) then hist448 <= hist448 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*449) and (unsigned(time_tmp) <= unsigned(delta)*450) ) then hist449 <= hist449 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*450) and (unsigned(time_tmp) <= unsigned(delta)*451) ) then hist450 <= hist450 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*451) and (unsigned(time_tmp) <= unsigned(delta)*452) ) then hist451 <= hist451 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*452) and (unsigned(time_tmp) <= unsigned(delta)*453) ) then hist452 <= hist452 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*453) and (unsigned(time_tmp) <= unsigned(delta)*454) ) then hist453 <= hist453 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*454) and (unsigned(time_tmp) <= unsigned(delta)*455) ) then hist454 <= hist454 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*455) and (unsigned(time_tmp) <= unsigned(delta)*456) ) then hist455 <= hist455 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*456) and (unsigned(time_tmp) <= unsigned(delta)*457) ) then hist456 <= hist456 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*457) and (unsigned(time_tmp) <= unsigned(delta)*458) ) then hist457 <= hist457 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*458) and (unsigned(time_tmp) <= unsigned(delta)*459) ) then hist458 <= hist458 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*459) and (unsigned(time_tmp) <= unsigned(delta)*460) ) then hist459 <= hist459 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*460) and (unsigned(time_tmp) <= unsigned(delta)*461) ) then hist460 <= hist460 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*461) and (unsigned(time_tmp) <= unsigned(delta)*462) ) then hist461 <= hist461 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*462) and (unsigned(time_tmp) <= unsigned(delta)*463) ) then hist462 <= hist462 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*463) and (unsigned(time_tmp) <= unsigned(delta)*464) ) then hist463 <= hist463 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*464) and (unsigned(time_tmp) <= unsigned(delta)*465) ) then hist464 <= hist464 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*465) and (unsigned(time_tmp) <= unsigned(delta)*466) ) then hist465 <= hist465 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*466) and (unsigned(time_tmp) <= unsigned(delta)*467) ) then hist466 <= hist466 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*467) and (unsigned(time_tmp) <= unsigned(delta)*468) ) then hist467 <= hist467 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*468) and (unsigned(time_tmp) <= unsigned(delta)*469) ) then hist468 <= hist468 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*469) and (unsigned(time_tmp) <= unsigned(delta)*470) ) then hist469 <= hist469 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*470) and (unsigned(time_tmp) <= unsigned(delta)*471) ) then hist470 <= hist470 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*471) and (unsigned(time_tmp) <= unsigned(delta)*472) ) then hist471 <= hist471 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*472) and (unsigned(time_tmp) <= unsigned(delta)*473) ) then hist472 <= hist472 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*473) and (unsigned(time_tmp) <= unsigned(delta)*474) ) then hist473 <= hist473 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*474) and (unsigned(time_tmp) <= unsigned(delta)*475) ) then hist474 <= hist474 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*475) and (unsigned(time_tmp) <= unsigned(delta)*476) ) then hist475 <= hist475 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*476) and (unsigned(time_tmp) <= unsigned(delta)*477) ) then hist476 <= hist476 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*477) and (unsigned(time_tmp) <= unsigned(delta)*478) ) then hist477 <= hist477 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*478) and (unsigned(time_tmp) <= unsigned(delta)*479) ) then hist478 <= hist478 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*479) and (unsigned(time_tmp) <= unsigned(delta)*480) ) then hist479 <= hist479 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*480) and (unsigned(time_tmp) <= unsigned(delta)*481) ) then hist480 <= hist480 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*481) and (unsigned(time_tmp) <= unsigned(delta)*482) ) then hist481 <= hist481 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*482) and (unsigned(time_tmp) <= unsigned(delta)*483) ) then hist482 <= hist482 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*483) and (unsigned(time_tmp) <= unsigned(delta)*484) ) then hist483 <= hist483 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*484) and (unsigned(time_tmp) <= unsigned(delta)*485) ) then hist484 <= hist484 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*485) and (unsigned(time_tmp) <= unsigned(delta)*486) ) then hist485 <= hist485 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*486) and (unsigned(time_tmp) <= unsigned(delta)*487) ) then hist486 <= hist486 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*487) and (unsigned(time_tmp) <= unsigned(delta)*488) ) then hist487 <= hist487 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*488) and (unsigned(time_tmp) <= unsigned(delta)*489) ) then hist488 <= hist488 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*489) and (unsigned(time_tmp) <= unsigned(delta)*490) ) then hist489 <= hist489 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*490) and (unsigned(time_tmp) <= unsigned(delta)*491) ) then hist490 <= hist490 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*491) and (unsigned(time_tmp) <= unsigned(delta)*492) ) then hist491 <= hist491 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*492) and (unsigned(time_tmp) <= unsigned(delta)*493) ) then hist492 <= hist492 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*493) and (unsigned(time_tmp) <= unsigned(delta)*494) ) then hist493 <= hist493 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*494) and (unsigned(time_tmp) <= unsigned(delta)*495) ) then hist494 <= hist494 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*495) and (unsigned(time_tmp) <= unsigned(delta)*496) ) then hist495 <= hist495 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*496) and (unsigned(time_tmp) <= unsigned(delta)*497) ) then hist496 <= hist496 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*497) and (unsigned(time_tmp) <= unsigned(delta)*498) ) then hist497 <= hist497 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*498) and (unsigned(time_tmp) <= unsigned(delta)*499) ) then hist498 <= hist498 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*499) and (unsigned(time_tmp) <= unsigned(delta)*500) ) then hist499 <= hist499 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*500) and (unsigned(time_tmp) <= unsigned(delta)*501) ) then hist500 <= hist500 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*501) and (unsigned(time_tmp) <= unsigned(delta)*502) ) then hist501 <= hist501 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*502) and (unsigned(time_tmp) <= unsigned(delta)*503) ) then hist502 <= hist502 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*503) and (unsigned(time_tmp) <= unsigned(delta)*504) ) then hist503 <= hist503 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*504) and (unsigned(time_tmp) <= unsigned(delta)*505) ) then hist504 <= hist504 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*505) and (unsigned(time_tmp) <= unsigned(delta)*506) ) then hist505 <= hist505 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*506) and (unsigned(time_tmp) <= unsigned(delta)*507) ) then hist506 <= hist506 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*507) and (unsigned(time_tmp) <= unsigned(delta)*508) ) then hist507 <= hist507 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*508) and (unsigned(time_tmp) <= unsigned(delta)*509) ) then hist508 <= hist508 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*509) and (unsigned(time_tmp) <= unsigned(delta)*510) ) then hist509 <= hist509 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*510) and (unsigned(time_tmp) <= unsigned(delta)*511) ) then hist510 <= hist510 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*511) and (unsigned(time_tmp) <= unsigned(delta)*512) ) then hist511 <= hist511 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*512) and (unsigned(time_tmp) <= unsigned(delta)*513) ) then hist512 <= hist512 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*513) and (unsigned(time_tmp) <= unsigned(delta)*514) ) then hist513 <= hist513 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*514) and (unsigned(time_tmp) <= unsigned(delta)*515) ) then hist514 <= hist514 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*515) and (unsigned(time_tmp) <= unsigned(delta)*516) ) then hist515 <= hist515 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*516) and (unsigned(time_tmp) <= unsigned(delta)*517) ) then hist516 <= hist516 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*517) and (unsigned(time_tmp) <= unsigned(delta)*518) ) then hist517 <= hist517 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*518) and (unsigned(time_tmp) <= unsigned(delta)*519) ) then hist518 <= hist518 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*519) and (unsigned(time_tmp) <= unsigned(delta)*520) ) then hist519 <= hist519 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*520) and (unsigned(time_tmp) <= unsigned(delta)*521) ) then hist520 <= hist520 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*521) and (unsigned(time_tmp) <= unsigned(delta)*522) ) then hist521 <= hist521 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*522) and (unsigned(time_tmp) <= unsigned(delta)*523) ) then hist522 <= hist522 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*523) and (unsigned(time_tmp) <= unsigned(delta)*524) ) then hist523 <= hist523 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*524) and (unsigned(time_tmp) <= unsigned(delta)*525) ) then hist524 <= hist524 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*525) and (unsigned(time_tmp) <= unsigned(delta)*526) ) then hist525 <= hist525 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*526) and (unsigned(time_tmp) <= unsigned(delta)*527) ) then hist526 <= hist526 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*527) and (unsigned(time_tmp) <= unsigned(delta)*528) ) then hist527 <= hist527 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*528) and (unsigned(time_tmp) <= unsigned(delta)*529) ) then hist528 <= hist528 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*529) and (unsigned(time_tmp) <= unsigned(delta)*530) ) then hist529 <= hist529 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*530) and (unsigned(time_tmp) <= unsigned(delta)*531) ) then hist530 <= hist530 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*531) and (unsigned(time_tmp) <= unsigned(delta)*532) ) then hist531 <= hist531 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*532) and (unsigned(time_tmp) <= unsigned(delta)*533) ) then hist532 <= hist532 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*533) and (unsigned(time_tmp) <= unsigned(delta)*534) ) then hist533 <= hist533 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*534) and (unsigned(time_tmp) <= unsigned(delta)*535) ) then hist534 <= hist534 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*535) and (unsigned(time_tmp) <= unsigned(delta)*536) ) then hist535 <= hist535 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*536) and (unsigned(time_tmp) <= unsigned(delta)*537) ) then hist536 <= hist536 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*537) and (unsigned(time_tmp) <= unsigned(delta)*538) ) then hist537 <= hist537 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*538) and (unsigned(time_tmp) <= unsigned(delta)*539) ) then hist538 <= hist538 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*539) and (unsigned(time_tmp) <= unsigned(delta)*540) ) then hist539 <= hist539 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*540) and (unsigned(time_tmp) <= unsigned(delta)*541) ) then hist540 <= hist540 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*541) and (unsigned(time_tmp) <= unsigned(delta)*542) ) then hist541 <= hist541 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*542) and (unsigned(time_tmp) <= unsigned(delta)*543) ) then hist542 <= hist542 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*543) and (unsigned(time_tmp) <= unsigned(delta)*544) ) then hist543 <= hist543 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*544) and (unsigned(time_tmp) <= unsigned(delta)*545) ) then hist544 <= hist544 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*545) and (unsigned(time_tmp) <= unsigned(delta)*546) ) then hist545 <= hist545 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*546) and (unsigned(time_tmp) <= unsigned(delta)*547) ) then hist546 <= hist546 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*547) and (unsigned(time_tmp) <= unsigned(delta)*548) ) then hist547 <= hist547 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*548) and (unsigned(time_tmp) <= unsigned(delta)*549) ) then hist548 <= hist548 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*549) and (unsigned(time_tmp) <= unsigned(delta)*550) ) then hist549 <= hist549 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*550) and (unsigned(time_tmp) <= unsigned(delta)*551) ) then hist550 <= hist550 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*551) and (unsigned(time_tmp) <= unsigned(delta)*552) ) then hist551 <= hist551 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*552) and (unsigned(time_tmp) <= unsigned(delta)*553) ) then hist552 <= hist552 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*553) and (unsigned(time_tmp) <= unsigned(delta)*554) ) then hist553 <= hist553 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*554) and (unsigned(time_tmp) <= unsigned(delta)*555) ) then hist554 <= hist554 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*555) and (unsigned(time_tmp) <= unsigned(delta)*556) ) then hist555 <= hist555 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*556) and (unsigned(time_tmp) <= unsigned(delta)*557) ) then hist556 <= hist556 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*557) and (unsigned(time_tmp) <= unsigned(delta)*558) ) then hist557 <= hist557 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*558) and (unsigned(time_tmp) <= unsigned(delta)*559) ) then hist558 <= hist558 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*559) and (unsigned(time_tmp) <= unsigned(delta)*560) ) then hist559 <= hist559 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*560) and (unsigned(time_tmp) <= unsigned(delta)*561) ) then hist560 <= hist560 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*561) and (unsigned(time_tmp) <= unsigned(delta)*562) ) then hist561 <= hist561 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*562) and (unsigned(time_tmp) <= unsigned(delta)*563) ) then hist562 <= hist562 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*563) and (unsigned(time_tmp) <= unsigned(delta)*564) ) then hist563 <= hist563 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*564) and (unsigned(time_tmp) <= unsigned(delta)*565) ) then hist564 <= hist564 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*565) and (unsigned(time_tmp) <= unsigned(delta)*566) ) then hist565 <= hist565 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*566) and (unsigned(time_tmp) <= unsigned(delta)*567) ) then hist566 <= hist566 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*567) and (unsigned(time_tmp) <= unsigned(delta)*568) ) then hist567 <= hist567 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*568) and (unsigned(time_tmp) <= unsigned(delta)*569) ) then hist568 <= hist568 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*569) and (unsigned(time_tmp) <= unsigned(delta)*570) ) then hist569 <= hist569 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*570) and (unsigned(time_tmp) <= unsigned(delta)*571) ) then hist570 <= hist570 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*571) and (unsigned(time_tmp) <= unsigned(delta)*572) ) then hist571 <= hist571 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*572) and (unsigned(time_tmp) <= unsigned(delta)*573) ) then hist572 <= hist572 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*573) and (unsigned(time_tmp) <= unsigned(delta)*574) ) then hist573 <= hist573 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*574) and (unsigned(time_tmp) <= unsigned(delta)*575) ) then hist574 <= hist574 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*575) and (unsigned(time_tmp) <= unsigned(delta)*576) ) then hist575 <= hist575 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*576) and (unsigned(time_tmp) <= unsigned(delta)*577) ) then hist576 <= hist576 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*577) and (unsigned(time_tmp) <= unsigned(delta)*578) ) then hist577 <= hist577 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*578) and (unsigned(time_tmp) <= unsigned(delta)*579) ) then hist578 <= hist578 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*579) and (unsigned(time_tmp) <= unsigned(delta)*580) ) then hist579 <= hist579 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*580) and (unsigned(time_tmp) <= unsigned(delta)*581) ) then hist580 <= hist580 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*581) and (unsigned(time_tmp) <= unsigned(delta)*582) ) then hist581 <= hist581 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*582) and (unsigned(time_tmp) <= unsigned(delta)*583) ) then hist582 <= hist582 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*583) and (unsigned(time_tmp) <= unsigned(delta)*584) ) then hist583 <= hist583 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*584) and (unsigned(time_tmp) <= unsigned(delta)*585) ) then hist584 <= hist584 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*585) and (unsigned(time_tmp) <= unsigned(delta)*586) ) then hist585 <= hist585 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*586) and (unsigned(time_tmp) <= unsigned(delta)*587) ) then hist586 <= hist586 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*587) and (unsigned(time_tmp) <= unsigned(delta)*588) ) then hist587 <= hist587 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*588) and (unsigned(time_tmp) <= unsigned(delta)*589) ) then hist588 <= hist588 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*589) and (unsigned(time_tmp) <= unsigned(delta)*590) ) then hist589 <= hist589 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*590) and (unsigned(time_tmp) <= unsigned(delta)*591) ) then hist590 <= hist590 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*591) and (unsigned(time_tmp) <= unsigned(delta)*592) ) then hist591 <= hist591 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*592) and (unsigned(time_tmp) <= unsigned(delta)*593) ) then hist592 <= hist592 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*593) and (unsigned(time_tmp) <= unsigned(delta)*594) ) then hist593 <= hist593 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*594) and (unsigned(time_tmp) <= unsigned(delta)*595) ) then hist594 <= hist594 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*595) and (unsigned(time_tmp) <= unsigned(delta)*596) ) then hist595 <= hist595 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*596) and (unsigned(time_tmp) <= unsigned(delta)*597) ) then hist596 <= hist596 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*597) and (unsigned(time_tmp) <= unsigned(delta)*598) ) then hist597 <= hist597 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*598) and (unsigned(time_tmp) <= unsigned(delta)*599) ) then hist598 <= hist598 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*599) and (unsigned(time_tmp) <= unsigned(delta)*600) ) then hist599 <= hist599 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*600) and (unsigned(time_tmp) <= unsigned(delta)*601) ) then hist600 <= hist600 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*601) and (unsigned(time_tmp) <= unsigned(delta)*602) ) then hist601 <= hist601 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*602) and (unsigned(time_tmp) <= unsigned(delta)*603) ) then hist602 <= hist602 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*603) and (unsigned(time_tmp) <= unsigned(delta)*604) ) then hist603 <= hist603 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*604) and (unsigned(time_tmp) <= unsigned(delta)*605) ) then hist604 <= hist604 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*605) and (unsigned(time_tmp) <= unsigned(delta)*606) ) then hist605 <= hist605 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*606) and (unsigned(time_tmp) <= unsigned(delta)*607) ) then hist606 <= hist606 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*607) and (unsigned(time_tmp) <= unsigned(delta)*608) ) then hist607 <= hist607 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*608) and (unsigned(time_tmp) <= unsigned(delta)*609) ) then hist608 <= hist608 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*609) and (unsigned(time_tmp) <= unsigned(delta)*610) ) then hist609 <= hist609 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*610) and (unsigned(time_tmp) <= unsigned(delta)*611) ) then hist610 <= hist610 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*611) and (unsigned(time_tmp) <= unsigned(delta)*612) ) then hist611 <= hist611 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*612) and (unsigned(time_tmp) <= unsigned(delta)*613) ) then hist612 <= hist612 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*613) and (unsigned(time_tmp) <= unsigned(delta)*614) ) then hist613 <= hist613 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*614) and (unsigned(time_tmp) <= unsigned(delta)*615) ) then hist614 <= hist614 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*615) and (unsigned(time_tmp) <= unsigned(delta)*616) ) then hist615 <= hist615 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*616) and (unsigned(time_tmp) <= unsigned(delta)*617) ) then hist616 <= hist616 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*617) and (unsigned(time_tmp) <= unsigned(delta)*618) ) then hist617 <= hist617 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*618) and (unsigned(time_tmp) <= unsigned(delta)*619) ) then hist618 <= hist618 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*619) and (unsigned(time_tmp) <= unsigned(delta)*620) ) then hist619 <= hist619 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*620) and (unsigned(time_tmp) <= unsigned(delta)*621) ) then hist620 <= hist620 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*621) and (unsigned(time_tmp) <= unsigned(delta)*622) ) then hist621 <= hist621 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*622) and (unsigned(time_tmp) <= unsigned(delta)*623) ) then hist622 <= hist622 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*623) and (unsigned(time_tmp) <= unsigned(delta)*624) ) then hist623 <= hist623 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*624) and (unsigned(time_tmp) <= unsigned(delta)*625) ) then hist624 <= hist624 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*625) and (unsigned(time_tmp) <= unsigned(delta)*626) ) then hist625 <= hist625 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*626) and (unsigned(time_tmp) <= unsigned(delta)*627) ) then hist626 <= hist626 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*627) and (unsigned(time_tmp) <= unsigned(delta)*628) ) then hist627 <= hist627 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*628) and (unsigned(time_tmp) <= unsigned(delta)*629) ) then hist628 <= hist628 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*629) and (unsigned(time_tmp) <= unsigned(delta)*630) ) then hist629 <= hist629 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*630) and (unsigned(time_tmp) <= unsigned(delta)*631) ) then hist630 <= hist630 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*631) and (unsigned(time_tmp) <= unsigned(delta)*632) ) then hist631 <= hist631 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*632) and (unsigned(time_tmp) <= unsigned(delta)*633) ) then hist632 <= hist632 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*633) and (unsigned(time_tmp) <= unsigned(delta)*634) ) then hist633 <= hist633 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*634) and (unsigned(time_tmp) <= unsigned(delta)*635) ) then hist634 <= hist634 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*635) and (unsigned(time_tmp) <= unsigned(delta)*636) ) then hist635 <= hist635 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*636) and (unsigned(time_tmp) <= unsigned(delta)*637) ) then hist636 <= hist636 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*637) and (unsigned(time_tmp) <= unsigned(delta)*638) ) then hist637 <= hist637 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*638) and (unsigned(time_tmp) <= unsigned(delta)*639) ) then hist638 <= hist638 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*639) and (unsigned(time_tmp) <= unsigned(delta)*640) ) then hist639 <= hist639 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*640) and (unsigned(time_tmp) <= unsigned(delta)*641) ) then hist640 <= hist640 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*641) and (unsigned(time_tmp) <= unsigned(delta)*642) ) then hist641 <= hist641 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*642) and (unsigned(time_tmp) <= unsigned(delta)*643) ) then hist642 <= hist642 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*643) and (unsigned(time_tmp) <= unsigned(delta)*644) ) then hist643 <= hist643 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*644) and (unsigned(time_tmp) <= unsigned(delta)*645) ) then hist644 <= hist644 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*645) and (unsigned(time_tmp) <= unsigned(delta)*646) ) then hist645 <= hist645 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*646) and (unsigned(time_tmp) <= unsigned(delta)*647) ) then hist646 <= hist646 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*647) and (unsigned(time_tmp) <= unsigned(delta)*648) ) then hist647 <= hist647 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*648) and (unsigned(time_tmp) <= unsigned(delta)*649) ) then hist648 <= hist648 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*649) and (unsigned(time_tmp) <= unsigned(delta)*650) ) then hist649 <= hist649 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*650) and (unsigned(time_tmp) <= unsigned(delta)*651) ) then hist650 <= hist650 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*651) and (unsigned(time_tmp) <= unsigned(delta)*652) ) then hist651 <= hist651 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*652) and (unsigned(time_tmp) <= unsigned(delta)*653) ) then hist652 <= hist652 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*653) and (unsigned(time_tmp) <= unsigned(delta)*654) ) then hist653 <= hist653 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*654) and (unsigned(time_tmp) <= unsigned(delta)*655) ) then hist654 <= hist654 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*655) and (unsigned(time_tmp) <= unsigned(delta)*656) ) then hist655 <= hist655 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*656) and (unsigned(time_tmp) <= unsigned(delta)*657) ) then hist656 <= hist656 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*657) and (unsigned(time_tmp) <= unsigned(delta)*658) ) then hist657 <= hist657 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*658) and (unsigned(time_tmp) <= unsigned(delta)*659) ) then hist658 <= hist658 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*659) and (unsigned(time_tmp) <= unsigned(delta)*660) ) then hist659 <= hist659 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*660) and (unsigned(time_tmp) <= unsigned(delta)*661) ) then hist660 <= hist660 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*661) and (unsigned(time_tmp) <= unsigned(delta)*662) ) then hist661 <= hist661 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*662) and (unsigned(time_tmp) <= unsigned(delta)*663) ) then hist662 <= hist662 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*663) and (unsigned(time_tmp) <= unsigned(delta)*664) ) then hist663 <= hist663 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*664) and (unsigned(time_tmp) <= unsigned(delta)*665) ) then hist664 <= hist664 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*665) and (unsigned(time_tmp) <= unsigned(delta)*666) ) then hist665 <= hist665 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*666) and (unsigned(time_tmp) <= unsigned(delta)*667) ) then hist666 <= hist666 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*667) and (unsigned(time_tmp) <= unsigned(delta)*668) ) then hist667 <= hist667 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*668) and (unsigned(time_tmp) <= unsigned(delta)*669) ) then hist668 <= hist668 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*669) and (unsigned(time_tmp) <= unsigned(delta)*670) ) then hist669 <= hist669 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*670) and (unsigned(time_tmp) <= unsigned(delta)*671) ) then hist670 <= hist670 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*671) and (unsigned(time_tmp) <= unsigned(delta)*672) ) then hist671 <= hist671 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*672) and (unsigned(time_tmp) <= unsigned(delta)*673) ) then hist672 <= hist672 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*673) and (unsigned(time_tmp) <= unsigned(delta)*674) ) then hist673 <= hist673 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*674) and (unsigned(time_tmp) <= unsigned(delta)*675) ) then hist674 <= hist674 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*675) and (unsigned(time_tmp) <= unsigned(delta)*676) ) then hist675 <= hist675 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*676) and (unsigned(time_tmp) <= unsigned(delta)*677) ) then hist676 <= hist676 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*677) and (unsigned(time_tmp) <= unsigned(delta)*678) ) then hist677 <= hist677 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*678) and (unsigned(time_tmp) <= unsigned(delta)*679) ) then hist678 <= hist678 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*679) and (unsigned(time_tmp) <= unsigned(delta)*680) ) then hist679 <= hist679 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*680) and (unsigned(time_tmp) <= unsigned(delta)*681) ) then hist680 <= hist680 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*681) and (unsigned(time_tmp) <= unsigned(delta)*682) ) then hist681 <= hist681 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*682) and (unsigned(time_tmp) <= unsigned(delta)*683) ) then hist682 <= hist682 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*683) and (unsigned(time_tmp) <= unsigned(delta)*684) ) then hist683 <= hist683 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*684) and (unsigned(time_tmp) <= unsigned(delta)*685) ) then hist684 <= hist684 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*685) and (unsigned(time_tmp) <= unsigned(delta)*686) ) then hist685 <= hist685 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*686) and (unsigned(time_tmp) <= unsigned(delta)*687) ) then hist686 <= hist686 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*687) and (unsigned(time_tmp) <= unsigned(delta)*688) ) then hist687 <= hist687 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*688) and (unsigned(time_tmp) <= unsigned(delta)*689) ) then hist688 <= hist688 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*689) and (unsigned(time_tmp) <= unsigned(delta)*690) ) then hist689 <= hist689 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*690) and (unsigned(time_tmp) <= unsigned(delta)*691) ) then hist690 <= hist690 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*691) and (unsigned(time_tmp) <= unsigned(delta)*692) ) then hist691 <= hist691 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*692) and (unsigned(time_tmp) <= unsigned(delta)*693) ) then hist692 <= hist692 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*693) and (unsigned(time_tmp) <= unsigned(delta)*694) ) then hist693 <= hist693 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*694) and (unsigned(time_tmp) <= unsigned(delta)*695) ) then hist694 <= hist694 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*695) and (unsigned(time_tmp) <= unsigned(delta)*696) ) then hist695 <= hist695 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*696) and (unsigned(time_tmp) <= unsigned(delta)*697) ) then hist696 <= hist696 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*697) and (unsigned(time_tmp) <= unsigned(delta)*698) ) then hist697 <= hist697 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*698) and (unsigned(time_tmp) <= unsigned(delta)*699) ) then hist698 <= hist698 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*699) and (unsigned(time_tmp) <= unsigned(delta)*700) ) then hist699 <= hist699 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*700) and (unsigned(time_tmp) <= unsigned(delta)*701) ) then hist700 <= hist700 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*701) and (unsigned(time_tmp) <= unsigned(delta)*702) ) then hist701 <= hist701 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*702) and (unsigned(time_tmp) <= unsigned(delta)*703) ) then hist702 <= hist702 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*703) and (unsigned(time_tmp) <= unsigned(delta)*704) ) then hist703 <= hist703 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*704) and (unsigned(time_tmp) <= unsigned(delta)*705) ) then hist704 <= hist704 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*705) and (unsigned(time_tmp) <= unsigned(delta)*706) ) then hist705 <= hist705 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*706) and (unsigned(time_tmp) <= unsigned(delta)*707) ) then hist706 <= hist706 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*707) and (unsigned(time_tmp) <= unsigned(delta)*708) ) then hist707 <= hist707 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*708) and (unsigned(time_tmp) <= unsigned(delta)*709) ) then hist708 <= hist708 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*709) and (unsigned(time_tmp) <= unsigned(delta)*710) ) then hist709 <= hist709 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*710) and (unsigned(time_tmp) <= unsigned(delta)*711) ) then hist710 <= hist710 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*711) and (unsigned(time_tmp) <= unsigned(delta)*712) ) then hist711 <= hist711 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*712) and (unsigned(time_tmp) <= unsigned(delta)*713) ) then hist712 <= hist712 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*713) and (unsigned(time_tmp) <= unsigned(delta)*714) ) then hist713 <= hist713 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*714) and (unsigned(time_tmp) <= unsigned(delta)*715) ) then hist714 <= hist714 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*715) and (unsigned(time_tmp) <= unsigned(delta)*716) ) then hist715 <= hist715 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*716) and (unsigned(time_tmp) <= unsigned(delta)*717) ) then hist716 <= hist716 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*717) and (unsigned(time_tmp) <= unsigned(delta)*718) ) then hist717 <= hist717 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*718) and (unsigned(time_tmp) <= unsigned(delta)*719) ) then hist718 <= hist718 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*719) and (unsigned(time_tmp) <= unsigned(delta)*720) ) then hist719 <= hist719 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*720) and (unsigned(time_tmp) <= unsigned(delta)*721) ) then hist720 <= hist720 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*721) and (unsigned(time_tmp) <= unsigned(delta)*722) ) then hist721 <= hist721 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*722) and (unsigned(time_tmp) <= unsigned(delta)*723) ) then hist722 <= hist722 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*723) and (unsigned(time_tmp) <= unsigned(delta)*724) ) then hist723 <= hist723 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*724) and (unsigned(time_tmp) <= unsigned(delta)*725) ) then hist724 <= hist724 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*725) and (unsigned(time_tmp) <= unsigned(delta)*726) ) then hist725 <= hist725 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*726) and (unsigned(time_tmp) <= unsigned(delta)*727) ) then hist726 <= hist726 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*727) and (unsigned(time_tmp) <= unsigned(delta)*728) ) then hist727 <= hist727 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*728) and (unsigned(time_tmp) <= unsigned(delta)*729) ) then hist728 <= hist728 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*729) and (unsigned(time_tmp) <= unsigned(delta)*730) ) then hist729 <= hist729 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*730) and (unsigned(time_tmp) <= unsigned(delta)*731) ) then hist730 <= hist730 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*731) and (unsigned(time_tmp) <= unsigned(delta)*732) ) then hist731 <= hist731 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*732) and (unsigned(time_tmp) <= unsigned(delta)*733) ) then hist732 <= hist732 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*733) and (unsigned(time_tmp) <= unsigned(delta)*734) ) then hist733 <= hist733 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*734) and (unsigned(time_tmp) <= unsigned(delta)*735) ) then hist734 <= hist734 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*735) and (unsigned(time_tmp) <= unsigned(delta)*736) ) then hist735 <= hist735 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*736) and (unsigned(time_tmp) <= unsigned(delta)*737) ) then hist736 <= hist736 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*737) and (unsigned(time_tmp) <= unsigned(delta)*738) ) then hist737 <= hist737 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*738) and (unsigned(time_tmp) <= unsigned(delta)*739) ) then hist738 <= hist738 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*739) and (unsigned(time_tmp) <= unsigned(delta)*740) ) then hist739 <= hist739 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*740) and (unsigned(time_tmp) <= unsigned(delta)*741) ) then hist740 <= hist740 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*741) and (unsigned(time_tmp) <= unsigned(delta)*742) ) then hist741 <= hist741 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*742) and (unsigned(time_tmp) <= unsigned(delta)*743) ) then hist742 <= hist742 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*743) and (unsigned(time_tmp) <= unsigned(delta)*744) ) then hist743 <= hist743 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*744) and (unsigned(time_tmp) <= unsigned(delta)*745) ) then hist744 <= hist744 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*745) and (unsigned(time_tmp) <= unsigned(delta)*746) ) then hist745 <= hist745 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*746) and (unsigned(time_tmp) <= unsigned(delta)*747) ) then hist746 <= hist746 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*747) and (unsigned(time_tmp) <= unsigned(delta)*748) ) then hist747 <= hist747 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*748) and (unsigned(time_tmp) <= unsigned(delta)*749) ) then hist748 <= hist748 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*749) and (unsigned(time_tmp) <= unsigned(delta)*750) ) then hist749 <= hist749 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*750) and (unsigned(time_tmp) <= unsigned(delta)*751) ) then hist750 <= hist750 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*751) and (unsigned(time_tmp) <= unsigned(delta)*752) ) then hist751 <= hist751 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*752) and (unsigned(time_tmp) <= unsigned(delta)*753) ) then hist752 <= hist752 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*753) and (unsigned(time_tmp) <= unsigned(delta)*754) ) then hist753 <= hist753 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*754) and (unsigned(time_tmp) <= unsigned(delta)*755) ) then hist754 <= hist754 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*755) and (unsigned(time_tmp) <= unsigned(delta)*756) ) then hist755 <= hist755 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*756) and (unsigned(time_tmp) <= unsigned(delta)*757) ) then hist756 <= hist756 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*757) and (unsigned(time_tmp) <= unsigned(delta)*758) ) then hist757 <= hist757 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*758) and (unsigned(time_tmp) <= unsigned(delta)*759) ) then hist758 <= hist758 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*759) and (unsigned(time_tmp) <= unsigned(delta)*760) ) then hist759 <= hist759 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*760) and (unsigned(time_tmp) <= unsigned(delta)*761) ) then hist760 <= hist760 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*761) and (unsigned(time_tmp) <= unsigned(delta)*762) ) then hist761 <= hist761 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*762) and (unsigned(time_tmp) <= unsigned(delta)*763) ) then hist762 <= hist762 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*763) and (unsigned(time_tmp) <= unsigned(delta)*764) ) then hist763 <= hist763 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*764) and (unsigned(time_tmp) <= unsigned(delta)*765) ) then hist764 <= hist764 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*765) and (unsigned(time_tmp) <= unsigned(delta)*766) ) then hist765 <= hist765 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*766) and (unsigned(time_tmp) <= unsigned(delta)*767) ) then hist766 <= hist766 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*767) and (unsigned(time_tmp) <= unsigned(delta)*768) ) then hist767 <= hist767 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*768) and (unsigned(time_tmp) <= unsigned(delta)*769) ) then hist768 <= hist768 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*769) and (unsigned(time_tmp) <= unsigned(delta)*770) ) then hist769 <= hist769 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*770) and (unsigned(time_tmp) <= unsigned(delta)*771) ) then hist770 <= hist770 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*771) and (unsigned(time_tmp) <= unsigned(delta)*772) ) then hist771 <= hist771 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*772) and (unsigned(time_tmp) <= unsigned(delta)*773) ) then hist772 <= hist772 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*773) and (unsigned(time_tmp) <= unsigned(delta)*774) ) then hist773 <= hist773 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*774) and (unsigned(time_tmp) <= unsigned(delta)*775) ) then hist774 <= hist774 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*775) and (unsigned(time_tmp) <= unsigned(delta)*776) ) then hist775 <= hist775 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*776) and (unsigned(time_tmp) <= unsigned(delta)*777) ) then hist776 <= hist776 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*777) and (unsigned(time_tmp) <= unsigned(delta)*778) ) then hist777 <= hist777 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*778) and (unsigned(time_tmp) <= unsigned(delta)*779) ) then hist778 <= hist778 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*779) and (unsigned(time_tmp) <= unsigned(delta)*780) ) then hist779 <= hist779 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*780) and (unsigned(time_tmp) <= unsigned(delta)*781) ) then hist780 <= hist780 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*781) and (unsigned(time_tmp) <= unsigned(delta)*782) ) then hist781 <= hist781 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*782) and (unsigned(time_tmp) <= unsigned(delta)*783) ) then hist782 <= hist782 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*783) and (unsigned(time_tmp) <= unsigned(delta)*784) ) then hist783 <= hist783 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*784) and (unsigned(time_tmp) <= unsigned(delta)*785) ) then hist784 <= hist784 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*785) and (unsigned(time_tmp) <= unsigned(delta)*786) ) then hist785 <= hist785 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*786) and (unsigned(time_tmp) <= unsigned(delta)*787) ) then hist786 <= hist786 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*787) and (unsigned(time_tmp) <= unsigned(delta)*788) ) then hist787 <= hist787 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*788) and (unsigned(time_tmp) <= unsigned(delta)*789) ) then hist788 <= hist788 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*789) and (unsigned(time_tmp) <= unsigned(delta)*790) ) then hist789 <= hist789 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*790) and (unsigned(time_tmp) <= unsigned(delta)*791) ) then hist790 <= hist790 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*791) and (unsigned(time_tmp) <= unsigned(delta)*792) ) then hist791 <= hist791 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*792) and (unsigned(time_tmp) <= unsigned(delta)*793) ) then hist792 <= hist792 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*793) and (unsigned(time_tmp) <= unsigned(delta)*794) ) then hist793 <= hist793 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*794) and (unsigned(time_tmp) <= unsigned(delta)*795) ) then hist794 <= hist794 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*795) and (unsigned(time_tmp) <= unsigned(delta)*796) ) then hist795 <= hist795 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*796) and (unsigned(time_tmp) <= unsigned(delta)*797) ) then hist796 <= hist796 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*797) and (unsigned(time_tmp) <= unsigned(delta)*798) ) then hist797 <= hist797 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*798) and (unsigned(time_tmp) <= unsigned(delta)*799) ) then hist798 <= hist798 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*799) and (unsigned(time_tmp) <= unsigned(delta)*800) ) then hist799 <= hist799 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*800) and (unsigned(time_tmp) <= unsigned(delta)*801) ) then hist800 <= hist800 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*801) and (unsigned(time_tmp) <= unsigned(delta)*802) ) then hist801 <= hist801 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*802) and (unsigned(time_tmp) <= unsigned(delta)*803) ) then hist802 <= hist802 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*803) and (unsigned(time_tmp) <= unsigned(delta)*804) ) then hist803 <= hist803 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*804) and (unsigned(time_tmp) <= unsigned(delta)*805) ) then hist804 <= hist804 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*805) and (unsigned(time_tmp) <= unsigned(delta)*806) ) then hist805 <= hist805 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*806) and (unsigned(time_tmp) <= unsigned(delta)*807) ) then hist806 <= hist806 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*807) and (unsigned(time_tmp) <= unsigned(delta)*808) ) then hist807 <= hist807 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*808) and (unsigned(time_tmp) <= unsigned(delta)*809) ) then hist808 <= hist808 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*809) and (unsigned(time_tmp) <= unsigned(delta)*810) ) then hist809 <= hist809 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*810) and (unsigned(time_tmp) <= unsigned(delta)*811) ) then hist810 <= hist810 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*811) and (unsigned(time_tmp) <= unsigned(delta)*812) ) then hist811 <= hist811 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*812) and (unsigned(time_tmp) <= unsigned(delta)*813) ) then hist812 <= hist812 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*813) and (unsigned(time_tmp) <= unsigned(delta)*814) ) then hist813 <= hist813 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*814) and (unsigned(time_tmp) <= unsigned(delta)*815) ) then hist814 <= hist814 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*815) and (unsigned(time_tmp) <= unsigned(delta)*816) ) then hist815 <= hist815 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*816) and (unsigned(time_tmp) <= unsigned(delta)*817) ) then hist816 <= hist816 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*817) and (unsigned(time_tmp) <= unsigned(delta)*818) ) then hist817 <= hist817 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*818) and (unsigned(time_tmp) <= unsigned(delta)*819) ) then hist818 <= hist818 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*819) and (unsigned(time_tmp) <= unsigned(delta)*820) ) then hist819 <= hist819 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*820) and (unsigned(time_tmp) <= unsigned(delta)*821) ) then hist820 <= hist820 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*821) and (unsigned(time_tmp) <= unsigned(delta)*822) ) then hist821 <= hist821 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*822) and (unsigned(time_tmp) <= unsigned(delta)*823) ) then hist822 <= hist822 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*823) and (unsigned(time_tmp) <= unsigned(delta)*824) ) then hist823 <= hist823 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*824) and (unsigned(time_tmp) <= unsigned(delta)*825) ) then hist824 <= hist824 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*825) and (unsigned(time_tmp) <= unsigned(delta)*826) ) then hist825 <= hist825 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*826) and (unsigned(time_tmp) <= unsigned(delta)*827) ) then hist826 <= hist826 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*827) and (unsigned(time_tmp) <= unsigned(delta)*828) ) then hist827 <= hist827 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*828) and (unsigned(time_tmp) <= unsigned(delta)*829) ) then hist828 <= hist828 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*829) and (unsigned(time_tmp) <= unsigned(delta)*830) ) then hist829 <= hist829 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*830) and (unsigned(time_tmp) <= unsigned(delta)*831) ) then hist830 <= hist830 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*831) and (unsigned(time_tmp) <= unsigned(delta)*832) ) then hist831 <= hist831 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*832) and (unsigned(time_tmp) <= unsigned(delta)*833) ) then hist832 <= hist832 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*833) and (unsigned(time_tmp) <= unsigned(delta)*834) ) then hist833 <= hist833 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*834) and (unsigned(time_tmp) <= unsigned(delta)*835) ) then hist834 <= hist834 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*835) and (unsigned(time_tmp) <= unsigned(delta)*836) ) then hist835 <= hist835 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*836) and (unsigned(time_tmp) <= unsigned(delta)*837) ) then hist836 <= hist836 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*837) and (unsigned(time_tmp) <= unsigned(delta)*838) ) then hist837 <= hist837 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*838) and (unsigned(time_tmp) <= unsigned(delta)*839) ) then hist838 <= hist838 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*839) and (unsigned(time_tmp) <= unsigned(delta)*840) ) then hist839 <= hist839 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*840) and (unsigned(time_tmp) <= unsigned(delta)*841) ) then hist840 <= hist840 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*841) and (unsigned(time_tmp) <= unsigned(delta)*842) ) then hist841 <= hist841 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*842) and (unsigned(time_tmp) <= unsigned(delta)*843) ) then hist842 <= hist842 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*843) and (unsigned(time_tmp) <= unsigned(delta)*844) ) then hist843 <= hist843 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*844) and (unsigned(time_tmp) <= unsigned(delta)*845) ) then hist844 <= hist844 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*845) and (unsigned(time_tmp) <= unsigned(delta)*846) ) then hist845 <= hist845 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*846) and (unsigned(time_tmp) <= unsigned(delta)*847) ) then hist846 <= hist846 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*847) and (unsigned(time_tmp) <= unsigned(delta)*848) ) then hist847 <= hist847 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*848) and (unsigned(time_tmp) <= unsigned(delta)*849) ) then hist848 <= hist848 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*849) and (unsigned(time_tmp) <= unsigned(delta)*850) ) then hist849 <= hist849 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*850) and (unsigned(time_tmp) <= unsigned(delta)*851) ) then hist850 <= hist850 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*851) and (unsigned(time_tmp) <= unsigned(delta)*852) ) then hist851 <= hist851 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*852) and (unsigned(time_tmp) <= unsigned(delta)*853) ) then hist852 <= hist852 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*853) and (unsigned(time_tmp) <= unsigned(delta)*854) ) then hist853 <= hist853 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*854) and (unsigned(time_tmp) <= unsigned(delta)*855) ) then hist854 <= hist854 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*855) and (unsigned(time_tmp) <= unsigned(delta)*856) ) then hist855 <= hist855 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*856) and (unsigned(time_tmp) <= unsigned(delta)*857) ) then hist856 <= hist856 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*857) and (unsigned(time_tmp) <= unsigned(delta)*858) ) then hist857 <= hist857 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*858) and (unsigned(time_tmp) <= unsigned(delta)*859) ) then hist858 <= hist858 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*859) and (unsigned(time_tmp) <= unsigned(delta)*860) ) then hist859 <= hist859 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*860) and (unsigned(time_tmp) <= unsigned(delta)*861) ) then hist860 <= hist860 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*861) and (unsigned(time_tmp) <= unsigned(delta)*862) ) then hist861 <= hist861 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*862) and (unsigned(time_tmp) <= unsigned(delta)*863) ) then hist862 <= hist862 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*863) and (unsigned(time_tmp) <= unsigned(delta)*864) ) then hist863 <= hist863 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*864) and (unsigned(time_tmp) <= unsigned(delta)*865) ) then hist864 <= hist864 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*865) and (unsigned(time_tmp) <= unsigned(delta)*866) ) then hist865 <= hist865 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*866) and (unsigned(time_tmp) <= unsigned(delta)*867) ) then hist866 <= hist866 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*867) and (unsigned(time_tmp) <= unsigned(delta)*868) ) then hist867 <= hist867 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*868) and (unsigned(time_tmp) <= unsigned(delta)*869) ) then hist868 <= hist868 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*869) and (unsigned(time_tmp) <= unsigned(delta)*870) ) then hist869 <= hist869 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*870) and (unsigned(time_tmp) <= unsigned(delta)*871) ) then hist870 <= hist870 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*871) and (unsigned(time_tmp) <= unsigned(delta)*872) ) then hist871 <= hist871 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*872) and (unsigned(time_tmp) <= unsigned(delta)*873) ) then hist872 <= hist872 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*873) and (unsigned(time_tmp) <= unsigned(delta)*874) ) then hist873 <= hist873 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*874) and (unsigned(time_tmp) <= unsigned(delta)*875) ) then hist874 <= hist874 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*875) and (unsigned(time_tmp) <= unsigned(delta)*876) ) then hist875 <= hist875 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*876) and (unsigned(time_tmp) <= unsigned(delta)*877) ) then hist876 <= hist876 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*877) and (unsigned(time_tmp) <= unsigned(delta)*878) ) then hist877 <= hist877 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*878) and (unsigned(time_tmp) <= unsigned(delta)*879) ) then hist878 <= hist878 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*879) and (unsigned(time_tmp) <= unsigned(delta)*880) ) then hist879 <= hist879 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*880) and (unsigned(time_tmp) <= unsigned(delta)*881) ) then hist880 <= hist880 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*881) and (unsigned(time_tmp) <= unsigned(delta)*882) ) then hist881 <= hist881 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*882) and (unsigned(time_tmp) <= unsigned(delta)*883) ) then hist882 <= hist882 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*883) and (unsigned(time_tmp) <= unsigned(delta)*884) ) then hist883 <= hist883 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*884) and (unsigned(time_tmp) <= unsigned(delta)*885) ) then hist884 <= hist884 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*885) and (unsigned(time_tmp) <= unsigned(delta)*886) ) then hist885 <= hist885 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*886) and (unsigned(time_tmp) <= unsigned(delta)*887) ) then hist886 <= hist886 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*887) and (unsigned(time_tmp) <= unsigned(delta)*888) ) then hist887 <= hist887 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*888) and (unsigned(time_tmp) <= unsigned(delta)*889) ) then hist888 <= hist888 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*889) and (unsigned(time_tmp) <= unsigned(delta)*890) ) then hist889 <= hist889 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*890) and (unsigned(time_tmp) <= unsigned(delta)*891) ) then hist890 <= hist890 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*891) and (unsigned(time_tmp) <= unsigned(delta)*892) ) then hist891 <= hist891 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*892) and (unsigned(time_tmp) <= unsigned(delta)*893) ) then hist892 <= hist892 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*893) and (unsigned(time_tmp) <= unsigned(delta)*894) ) then hist893 <= hist893 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*894) and (unsigned(time_tmp) <= unsigned(delta)*895) ) then hist894 <= hist894 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*895) and (unsigned(time_tmp) <= unsigned(delta)*896) ) then hist895 <= hist895 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*896) and (unsigned(time_tmp) <= unsigned(delta)*897) ) then hist896 <= hist896 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*897) and (unsigned(time_tmp) <= unsigned(delta)*898) ) then hist897 <= hist897 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*898) and (unsigned(time_tmp) <= unsigned(delta)*899) ) then hist898 <= hist898 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*899) and (unsigned(time_tmp) <= unsigned(delta)*900) ) then hist899 <= hist899 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*900) and (unsigned(time_tmp) <= unsigned(delta)*901) ) then hist900 <= hist900 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*901) and (unsigned(time_tmp) <= unsigned(delta)*902) ) then hist901 <= hist901 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*902) and (unsigned(time_tmp) <= unsigned(delta)*903) ) then hist902 <= hist902 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*903) and (unsigned(time_tmp) <= unsigned(delta)*904) ) then hist903 <= hist903 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*904) and (unsigned(time_tmp) <= unsigned(delta)*905) ) then hist904 <= hist904 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*905) and (unsigned(time_tmp) <= unsigned(delta)*906) ) then hist905 <= hist905 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*906) and (unsigned(time_tmp) <= unsigned(delta)*907) ) then hist906 <= hist906 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*907) and (unsigned(time_tmp) <= unsigned(delta)*908) ) then hist907 <= hist907 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*908) and (unsigned(time_tmp) <= unsigned(delta)*909) ) then hist908 <= hist908 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*909) and (unsigned(time_tmp) <= unsigned(delta)*910) ) then hist909 <= hist909 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*910) and (unsigned(time_tmp) <= unsigned(delta)*911) ) then hist910 <= hist910 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*911) and (unsigned(time_tmp) <= unsigned(delta)*912) ) then hist911 <= hist911 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*912) and (unsigned(time_tmp) <= unsigned(delta)*913) ) then hist912 <= hist912 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*913) and (unsigned(time_tmp) <= unsigned(delta)*914) ) then hist913 <= hist913 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*914) and (unsigned(time_tmp) <= unsigned(delta)*915) ) then hist914 <= hist914 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*915) and (unsigned(time_tmp) <= unsigned(delta)*916) ) then hist915 <= hist915 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*916) and (unsigned(time_tmp) <= unsigned(delta)*917) ) then hist916 <= hist916 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*917) and (unsigned(time_tmp) <= unsigned(delta)*918) ) then hist917 <= hist917 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*918) and (unsigned(time_tmp) <= unsigned(delta)*919) ) then hist918 <= hist918 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*919) and (unsigned(time_tmp) <= unsigned(delta)*920) ) then hist919 <= hist919 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*920) and (unsigned(time_tmp) <= unsigned(delta)*921) ) then hist920 <= hist920 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*921) and (unsigned(time_tmp) <= unsigned(delta)*922) ) then hist921 <= hist921 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*922) and (unsigned(time_tmp) <= unsigned(delta)*923) ) then hist922 <= hist922 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*923) and (unsigned(time_tmp) <= unsigned(delta)*924) ) then hist923 <= hist923 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*924) and (unsigned(time_tmp) <= unsigned(delta)*925) ) then hist924 <= hist924 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*925) and (unsigned(time_tmp) <= unsigned(delta)*926) ) then hist925 <= hist925 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*926) and (unsigned(time_tmp) <= unsigned(delta)*927) ) then hist926 <= hist926 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*927) and (unsigned(time_tmp) <= unsigned(delta)*928) ) then hist927 <= hist927 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*928) and (unsigned(time_tmp) <= unsigned(delta)*929) ) then hist928 <= hist928 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*929) and (unsigned(time_tmp) <= unsigned(delta)*930) ) then hist929 <= hist929 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*930) and (unsigned(time_tmp) <= unsigned(delta)*931) ) then hist930 <= hist930 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*931) and (unsigned(time_tmp) <= unsigned(delta)*932) ) then hist931 <= hist931 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*932) and (unsigned(time_tmp) <= unsigned(delta)*933) ) then hist932 <= hist932 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*933) and (unsigned(time_tmp) <= unsigned(delta)*934) ) then hist933 <= hist933 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*934) and (unsigned(time_tmp) <= unsigned(delta)*935) ) then hist934 <= hist934 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*935) and (unsigned(time_tmp) <= unsigned(delta)*936) ) then hist935 <= hist935 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*936) and (unsigned(time_tmp) <= unsigned(delta)*937) ) then hist936 <= hist936 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*937) and (unsigned(time_tmp) <= unsigned(delta)*938) ) then hist937 <= hist937 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*938) and (unsigned(time_tmp) <= unsigned(delta)*939) ) then hist938 <= hist938 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*939) and (unsigned(time_tmp) <= unsigned(delta)*940) ) then hist939 <= hist939 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*940) and (unsigned(time_tmp) <= unsigned(delta)*941) ) then hist940 <= hist940 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*941) and (unsigned(time_tmp) <= unsigned(delta)*942) ) then hist941 <= hist941 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*942) and (unsigned(time_tmp) <= unsigned(delta)*943) ) then hist942 <= hist942 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*943) and (unsigned(time_tmp) <= unsigned(delta)*944) ) then hist943 <= hist943 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*944) and (unsigned(time_tmp) <= unsigned(delta)*945) ) then hist944 <= hist944 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*945) and (unsigned(time_tmp) <= unsigned(delta)*946) ) then hist945 <= hist945 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*946) and (unsigned(time_tmp) <= unsigned(delta)*947) ) then hist946 <= hist946 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*947) and (unsigned(time_tmp) <= unsigned(delta)*948) ) then hist947 <= hist947 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*948) and (unsigned(time_tmp) <= unsigned(delta)*949) ) then hist948 <= hist948 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*949) and (unsigned(time_tmp) <= unsigned(delta)*950) ) then hist949 <= hist949 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*950) and (unsigned(time_tmp) <= unsigned(delta)*951) ) then hist950 <= hist950 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*951) and (unsigned(time_tmp) <= unsigned(delta)*952) ) then hist951 <= hist951 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*952) and (unsigned(time_tmp) <= unsigned(delta)*953) ) then hist952 <= hist952 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*953) and (unsigned(time_tmp) <= unsigned(delta)*954) ) then hist953 <= hist953 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*954) and (unsigned(time_tmp) <= unsigned(delta)*955) ) then hist954 <= hist954 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*955) and (unsigned(time_tmp) <= unsigned(delta)*956) ) then hist955 <= hist955 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*956) and (unsigned(time_tmp) <= unsigned(delta)*957) ) then hist956 <= hist956 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*957) and (unsigned(time_tmp) <= unsigned(delta)*958) ) then hist957 <= hist957 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*958) and (unsigned(time_tmp) <= unsigned(delta)*959) ) then hist958 <= hist958 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*959) and (unsigned(time_tmp) <= unsigned(delta)*960) ) then hist959 <= hist959 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*960) and (unsigned(time_tmp) <= unsigned(delta)*961) ) then hist960 <= hist960 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*961) and (unsigned(time_tmp) <= unsigned(delta)*962) ) then hist961 <= hist961 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*962) and (unsigned(time_tmp) <= unsigned(delta)*963) ) then hist962 <= hist962 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*963) and (unsigned(time_tmp) <= unsigned(delta)*964) ) then hist963 <= hist963 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*964) and (unsigned(time_tmp) <= unsigned(delta)*965) ) then hist964 <= hist964 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*965) and (unsigned(time_tmp) <= unsigned(delta)*966) ) then hist965 <= hist965 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*966) and (unsigned(time_tmp) <= unsigned(delta)*967) ) then hist966 <= hist966 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*967) and (unsigned(time_tmp) <= unsigned(delta)*968) ) then hist967 <= hist967 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*968) and (unsigned(time_tmp) <= unsigned(delta)*969) ) then hist968 <= hist968 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*969) and (unsigned(time_tmp) <= unsigned(delta)*970) ) then hist969 <= hist969 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*970) and (unsigned(time_tmp) <= unsigned(delta)*971) ) then hist970 <= hist970 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*971) and (unsigned(time_tmp) <= unsigned(delta)*972) ) then hist971 <= hist971 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*972) and (unsigned(time_tmp) <= unsigned(delta)*973) ) then hist972 <= hist972 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*973) and (unsigned(time_tmp) <= unsigned(delta)*974) ) then hist973 <= hist973 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*974) and (unsigned(time_tmp) <= unsigned(delta)*975) ) then hist974 <= hist974 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*975) and (unsigned(time_tmp) <= unsigned(delta)*976) ) then hist975 <= hist975 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*976) and (unsigned(time_tmp) <= unsigned(delta)*977) ) then hist976 <= hist976 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*977) and (unsigned(time_tmp) <= unsigned(delta)*978) ) then hist977 <= hist977 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*978) and (unsigned(time_tmp) <= unsigned(delta)*979) ) then hist978 <= hist978 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*979) and (unsigned(time_tmp) <= unsigned(delta)*980) ) then hist979 <= hist979 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*980) and (unsigned(time_tmp) <= unsigned(delta)*981) ) then hist980 <= hist980 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*981) and (unsigned(time_tmp) <= unsigned(delta)*982) ) then hist981 <= hist981 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*982) and (unsigned(time_tmp) <= unsigned(delta)*983) ) then hist982 <= hist982 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*983) and (unsigned(time_tmp) <= unsigned(delta)*984) ) then hist983 <= hist983 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*984) and (unsigned(time_tmp) <= unsigned(delta)*985) ) then hist984 <= hist984 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*985) and (unsigned(time_tmp) <= unsigned(delta)*986) ) then hist985 <= hist985 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*986) and (unsigned(time_tmp) <= unsigned(delta)*987) ) then hist986 <= hist986 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*987) and (unsigned(time_tmp) <= unsigned(delta)*988) ) then hist987 <= hist987 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*988) and (unsigned(time_tmp) <= unsigned(delta)*989) ) then hist988 <= hist988 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*989) and (unsigned(time_tmp) <= unsigned(delta)*990) ) then hist989 <= hist989 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*990) and (unsigned(time_tmp) <= unsigned(delta)*991) ) then hist990 <= hist990 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*991) and (unsigned(time_tmp) <= unsigned(delta)*992) ) then hist991 <= hist991 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*992) and (unsigned(time_tmp) <= unsigned(delta)*993) ) then hist992 <= hist992 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*993) and (unsigned(time_tmp) <= unsigned(delta)*994) ) then hist993 <= hist993 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*994) and (unsigned(time_tmp) <= unsigned(delta)*995) ) then hist994 <= hist994 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*995) and (unsigned(time_tmp) <= unsigned(delta)*996) ) then hist995 <= hist995 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*996) and (unsigned(time_tmp) <= unsigned(delta)*997) ) then hist996 <= hist996 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*997) and (unsigned(time_tmp) <= unsigned(delta)*998) ) then hist997 <= hist997 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*998) and (unsigned(time_tmp) <= unsigned(delta)*999) ) then hist998 <= hist998 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*999) and (unsigned(time_tmp) <= unsigned(delta)*1000) ) then hist999 <= hist999 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1000) and (unsigned(time_tmp) <= unsigned(delta)*1001) ) then hist1000 <= hist1000 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1001) and (unsigned(time_tmp) <= unsigned(delta)*1002) ) then hist1001 <= hist1001 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1002) and (unsigned(time_tmp) <= unsigned(delta)*1003) ) then hist1002 <= hist1002 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1003) and (unsigned(time_tmp) <= unsigned(delta)*1004) ) then hist1003 <= hist1003 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1004) and (unsigned(time_tmp) <= unsigned(delta)*1005) ) then hist1004 <= hist1004 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1005) and (unsigned(time_tmp) <= unsigned(delta)*1006) ) then hist1005 <= hist1005 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1006) and (unsigned(time_tmp) <= unsigned(delta)*1007) ) then hist1006 <= hist1006 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1007) and (unsigned(time_tmp) <= unsigned(delta)*1008) ) then hist1007 <= hist1007 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1008) and (unsigned(time_tmp) <= unsigned(delta)*1009) ) then hist1008 <= hist1008 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1009) and (unsigned(time_tmp) <= unsigned(delta)*1010) ) then hist1009 <= hist1009 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1010) and (unsigned(time_tmp) <= unsigned(delta)*1011) ) then hist1010 <= hist1010 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1011) and (unsigned(time_tmp) <= unsigned(delta)*1012) ) then hist1011 <= hist1011 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1012) and (unsigned(time_tmp) <= unsigned(delta)*1013) ) then hist1012 <= hist1012 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1013) and (unsigned(time_tmp) <= unsigned(delta)*1014) ) then hist1013 <= hist1013 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1014) and (unsigned(time_tmp) <= unsigned(delta)*1015) ) then hist1014 <= hist1014 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1015) and (unsigned(time_tmp) <= unsigned(delta)*1016) ) then hist1015 <= hist1015 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1016) and (unsigned(time_tmp) <= unsigned(delta)*1017) ) then hist1016 <= hist1016 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1017) and (unsigned(time_tmp) <= unsigned(delta)*1018) ) then hist1017 <= hist1017 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1018) and (unsigned(time_tmp) <= unsigned(delta)*1019) ) then hist1018 <= hist1018 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1019) and (unsigned(time_tmp) <= unsigned(delta)*1020) ) then hist1019 <= hist1019 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1020) and (unsigned(time_tmp) <= unsigned(delta)*1021) ) then hist1020 <= hist1020 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1021) and (unsigned(time_tmp) <= unsigned(delta)*1022) ) then hist1021 <= hist1021 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1022) and (unsigned(time_tmp) <= unsigned(delta)*1023) ) then hist1022 <= hist1022 + '1';
			elsif ((unsigned(time_tmp) > unsigned(delta)*1023) and (unsigned(time_tmp) <= unsigned(delta)*1024) ) then hist1023 <= hist1023 + '1';
			
			else

			end if;
	end if;	
	end if;	
	
end process;

--
hist( 31 downto 0 ) <= hist0 ( 31 downto 0 );
hist( 63 downto 32 ) <= hist1 ( 31 downto 0 );
hist( 95 downto 64 ) <= hist2 ( 31 downto 0 );
hist( 127 downto 96 ) <= hist3 ( 31 downto 0 );
hist( 159 downto 128 ) <= hist4 ( 31 downto 0 );
hist( 191 downto 160 ) <= hist5 ( 31 downto 0 );
hist( 223 downto 192 ) <= hist6 ( 31 downto 0 );
hist( 255 downto 224 ) <= hist7 ( 31 downto 0 );
hist( 287 downto 256 ) <= hist8 ( 31 downto 0 );
hist( 319 downto 288 ) <= hist9 ( 31 downto 0 );
hist( 351 downto 320 ) <= hist10 ( 31 downto 0 );
hist( 383 downto 352 ) <= hist11 ( 31 downto 0 );
hist( 415 downto 384 ) <= hist12 ( 31 downto 0 );
hist( 447 downto 416 ) <= hist13 ( 31 downto 0 );
hist( 479 downto 448 ) <= hist14 ( 31 downto 0 );
hist( 511 downto 480 ) <= hist15 ( 31 downto 0 );
hist( 543 downto 512 ) <= hist16 ( 31 downto 0 );
hist( 575 downto 544 ) <= hist17 ( 31 downto 0 );
hist( 607 downto 576 ) <= hist18 ( 31 downto 0 );
hist( 639 downto 608 ) <= hist19 ( 31 downto 0 );
hist( 671 downto 640 ) <= hist20 ( 31 downto 0 );
hist( 703 downto 672 ) <= hist21 ( 31 downto 0 );
hist( 735 downto 704 ) <= hist22 ( 31 downto 0 );
hist( 767 downto 736 ) <= hist23 ( 31 downto 0 );
hist( 799 downto 768 ) <= hist24 ( 31 downto 0 );
hist( 831 downto 800 ) <= hist25 ( 31 downto 0 );
hist( 863 downto 832 ) <= hist26 ( 31 downto 0 );
hist( 895 downto 864 ) <= hist27 ( 31 downto 0 );
hist( 927 downto 896 ) <= hist28 ( 31 downto 0 );
hist( 959 downto 928 ) <= hist29 ( 31 downto 0 );
hist( 991 downto 960 ) <= hist30 ( 31 downto 0 );
hist( 1023 downto 992 ) <= hist31 ( 31 downto 0 );
hist( 1055 downto 1024 ) <= hist32 ( 31 downto 0 );
hist( 1087 downto 1056 ) <= hist33 ( 31 downto 0 );
hist( 1119 downto 1088 ) <= hist34 ( 31 downto 0 );
hist( 1151 downto 1120 ) <= hist35 ( 31 downto 0 );
hist( 1183 downto 1152 ) <= hist36 ( 31 downto 0 );
hist( 1215 downto 1184 ) <= hist37 ( 31 downto 0 );
hist( 1247 downto 1216 ) <= hist38 ( 31 downto 0 );
hist( 1279 downto 1248 ) <= hist39 ( 31 downto 0 );
hist( 1311 downto 1280 ) <= hist40 ( 31 downto 0 );
hist( 1343 downto 1312 ) <= hist41 ( 31 downto 0 );
hist( 1375 downto 1344 ) <= hist42 ( 31 downto 0 );
hist( 1407 downto 1376 ) <= hist43 ( 31 downto 0 );
hist( 1439 downto 1408 ) <= hist44 ( 31 downto 0 );
hist( 1471 downto 1440 ) <= hist45 ( 31 downto 0 );
hist( 1503 downto 1472 ) <= hist46 ( 31 downto 0 );
hist( 1535 downto 1504 ) <= hist47 ( 31 downto 0 );
hist( 1567 downto 1536 ) <= hist48 ( 31 downto 0 );
hist( 1599 downto 1568 ) <= hist49 ( 31 downto 0 );
hist( 1631 downto 1600 ) <= hist50 ( 31 downto 0 );
hist( 1663 downto 1632 ) <= hist51 ( 31 downto 0 );
hist( 1695 downto 1664 ) <= hist52 ( 31 downto 0 );
hist( 1727 downto 1696 ) <= hist53 ( 31 downto 0 );
hist( 1759 downto 1728 ) <= hist54 ( 31 downto 0 );
hist( 1791 downto 1760 ) <= hist55 ( 31 downto 0 );
hist( 1823 downto 1792 ) <= hist56 ( 31 downto 0 );
hist( 1855 downto 1824 ) <= hist57 ( 31 downto 0 );
hist( 1887 downto 1856 ) <= hist58 ( 31 downto 0 );
hist( 1919 downto 1888 ) <= hist59 ( 31 downto 0 );
hist( 1951 downto 1920 ) <= hist60 ( 31 downto 0 );
hist( 1983 downto 1952 ) <= hist61 ( 31 downto 0 );
hist( 2015 downto 1984 ) <= hist62 ( 31 downto 0 );
hist( 2047 downto 2016 ) <= hist63 ( 31 downto 0 );
hist( 2079 downto 2048 ) <= hist64 ( 31 downto 0 );
hist( 2111 downto 2080 ) <= hist65 ( 31 downto 0 );
hist( 2143 downto 2112 ) <= hist66 ( 31 downto 0 );
hist( 2175 downto 2144 ) <= hist67 ( 31 downto 0 );
hist( 2207 downto 2176 ) <= hist68 ( 31 downto 0 );
hist( 2239 downto 2208 ) <= hist69 ( 31 downto 0 );
hist( 2271 downto 2240 ) <= hist70 ( 31 downto 0 );
hist( 2303 downto 2272 ) <= hist71 ( 31 downto 0 );
hist( 2335 downto 2304 ) <= hist72 ( 31 downto 0 );
hist( 2367 downto 2336 ) <= hist73 ( 31 downto 0 );
hist( 2399 downto 2368 ) <= hist74 ( 31 downto 0 );
hist( 2431 downto 2400 ) <= hist75 ( 31 downto 0 );
hist( 2463 downto 2432 ) <= hist76 ( 31 downto 0 );
hist( 2495 downto 2464 ) <= hist77 ( 31 downto 0 );
hist( 2527 downto 2496 ) <= hist78 ( 31 downto 0 );
hist( 2559 downto 2528 ) <= hist79 ( 31 downto 0 );
hist( 2591 downto 2560 ) <= hist80 ( 31 downto 0 );
hist( 2623 downto 2592 ) <= hist81 ( 31 downto 0 );
hist( 2655 downto 2624 ) <= hist82 ( 31 downto 0 );
hist( 2687 downto 2656 ) <= hist83 ( 31 downto 0 );
hist( 2719 downto 2688 ) <= hist84 ( 31 downto 0 );
hist( 2751 downto 2720 ) <= hist85 ( 31 downto 0 );
hist( 2783 downto 2752 ) <= hist86 ( 31 downto 0 );
hist( 2815 downto 2784 ) <= hist87 ( 31 downto 0 );
hist( 2847 downto 2816 ) <= hist88 ( 31 downto 0 );
hist( 2879 downto 2848 ) <= hist89 ( 31 downto 0 );
hist( 2911 downto 2880 ) <= hist90 ( 31 downto 0 );
hist( 2943 downto 2912 ) <= hist91 ( 31 downto 0 );
hist( 2975 downto 2944 ) <= hist92 ( 31 downto 0 );
hist( 3007 downto 2976 ) <= hist93 ( 31 downto 0 );
hist( 3039 downto 3008 ) <= hist94 ( 31 downto 0 );
hist( 3071 downto 3040 ) <= hist95 ( 31 downto 0 );
hist( 3103 downto 3072 ) <= hist96 ( 31 downto 0 );
hist( 3135 downto 3104 ) <= hist97 ( 31 downto 0 );
hist( 3167 downto 3136 ) <= hist98 ( 31 downto 0 );
hist( 3199 downto 3168 ) <= hist99 ( 31 downto 0 );
hist( 3231 downto 3200 ) <= hist100 ( 31 downto 0 );
hist( 3263 downto 3232 ) <= hist101 ( 31 downto 0 );
hist( 3295 downto 3264 ) <= hist102 ( 31 downto 0 );
hist( 3327 downto 3296 ) <= hist103 ( 31 downto 0 );
hist( 3359 downto 3328 ) <= hist104 ( 31 downto 0 );
hist( 3391 downto 3360 ) <= hist105 ( 31 downto 0 );
hist( 3423 downto 3392 ) <= hist106 ( 31 downto 0 );
hist( 3455 downto 3424 ) <= hist107 ( 31 downto 0 );
hist( 3487 downto 3456 ) <= hist108 ( 31 downto 0 );
hist( 3519 downto 3488 ) <= hist109 ( 31 downto 0 );
hist( 3551 downto 3520 ) <= hist110 ( 31 downto 0 );
hist( 3583 downto 3552 ) <= hist111 ( 31 downto 0 );
hist( 3615 downto 3584 ) <= hist112 ( 31 downto 0 );
hist( 3647 downto 3616 ) <= hist113 ( 31 downto 0 );
hist( 3679 downto 3648 ) <= hist114 ( 31 downto 0 );
hist( 3711 downto 3680 ) <= hist115 ( 31 downto 0 );
hist( 3743 downto 3712 ) <= hist116 ( 31 downto 0 );
hist( 3775 downto 3744 ) <= hist117 ( 31 downto 0 );
hist( 3807 downto 3776 ) <= hist118 ( 31 downto 0 );
hist( 3839 downto 3808 ) <= hist119 ( 31 downto 0 );
hist( 3871 downto 3840 ) <= hist120 ( 31 downto 0 );
hist( 3903 downto 3872 ) <= hist121 ( 31 downto 0 );
hist( 3935 downto 3904 ) <= hist122 ( 31 downto 0 );
hist( 3967 downto 3936 ) <= hist123 ( 31 downto 0 );
hist( 3999 downto 3968 ) <= hist124 ( 31 downto 0 );
hist( 4031 downto 4000 ) <= hist125 ( 31 downto 0 );
hist( 4063 downto 4032 ) <= hist126 ( 31 downto 0 );
hist( 4095 downto 4064 ) <= hist127 ( 31 downto 0 );
hist( 4127 downto 4096 ) <= hist128 ( 31 downto 0 );
hist( 4159 downto 4128 ) <= hist129 ( 31 downto 0 );
hist( 4191 downto 4160 ) <= hist130 ( 31 downto 0 );
hist( 4223 downto 4192 ) <= hist131 ( 31 downto 0 );
hist( 4255 downto 4224 ) <= hist132 ( 31 downto 0 );
hist( 4287 downto 4256 ) <= hist133 ( 31 downto 0 );
hist( 4319 downto 4288 ) <= hist134 ( 31 downto 0 );
hist( 4351 downto 4320 ) <= hist135 ( 31 downto 0 );
hist( 4383 downto 4352 ) <= hist136 ( 31 downto 0 );
hist( 4415 downto 4384 ) <= hist137 ( 31 downto 0 );
hist( 4447 downto 4416 ) <= hist138 ( 31 downto 0 );
hist( 4479 downto 4448 ) <= hist139 ( 31 downto 0 );
hist( 4511 downto 4480 ) <= hist140 ( 31 downto 0 );
hist( 4543 downto 4512 ) <= hist141 ( 31 downto 0 );
hist( 4575 downto 4544 ) <= hist142 ( 31 downto 0 );
hist( 4607 downto 4576 ) <= hist143 ( 31 downto 0 );
hist( 4639 downto 4608 ) <= hist144 ( 31 downto 0 );
hist( 4671 downto 4640 ) <= hist145 ( 31 downto 0 );
hist( 4703 downto 4672 ) <= hist146 ( 31 downto 0 );
hist( 4735 downto 4704 ) <= hist147 ( 31 downto 0 );
hist( 4767 downto 4736 ) <= hist148 ( 31 downto 0 );
hist( 4799 downto 4768 ) <= hist149 ( 31 downto 0 );
hist( 4831 downto 4800 ) <= hist150 ( 31 downto 0 );
hist( 4863 downto 4832 ) <= hist151 ( 31 downto 0 );
hist( 4895 downto 4864 ) <= hist152 ( 31 downto 0 );
hist( 4927 downto 4896 ) <= hist153 ( 31 downto 0 );
hist( 4959 downto 4928 ) <= hist154 ( 31 downto 0 );
hist( 4991 downto 4960 ) <= hist155 ( 31 downto 0 );
hist( 5023 downto 4992 ) <= hist156 ( 31 downto 0 );
hist( 5055 downto 5024 ) <= hist157 ( 31 downto 0 );
hist( 5087 downto 5056 ) <= hist158 ( 31 downto 0 );
hist( 5119 downto 5088 ) <= hist159 ( 31 downto 0 );
hist( 5151 downto 5120 ) <= hist160 ( 31 downto 0 );
hist( 5183 downto 5152 ) <= hist161 ( 31 downto 0 );
hist( 5215 downto 5184 ) <= hist162 ( 31 downto 0 );
hist( 5247 downto 5216 ) <= hist163 ( 31 downto 0 );
hist( 5279 downto 5248 ) <= hist164 ( 31 downto 0 );
hist( 5311 downto 5280 ) <= hist165 ( 31 downto 0 );
hist( 5343 downto 5312 ) <= hist166 ( 31 downto 0 );
hist( 5375 downto 5344 ) <= hist167 ( 31 downto 0 );
hist( 5407 downto 5376 ) <= hist168 ( 31 downto 0 );
hist( 5439 downto 5408 ) <= hist169 ( 31 downto 0 );
hist( 5471 downto 5440 ) <= hist170 ( 31 downto 0 );
hist( 5503 downto 5472 ) <= hist171 ( 31 downto 0 );
hist( 5535 downto 5504 ) <= hist172 ( 31 downto 0 );
hist( 5567 downto 5536 ) <= hist173 ( 31 downto 0 );
hist( 5599 downto 5568 ) <= hist174 ( 31 downto 0 );
hist( 5631 downto 5600 ) <= hist175 ( 31 downto 0 );
hist( 5663 downto 5632 ) <= hist176 ( 31 downto 0 );
hist( 5695 downto 5664 ) <= hist177 ( 31 downto 0 );
hist( 5727 downto 5696 ) <= hist178 ( 31 downto 0 );
hist( 5759 downto 5728 ) <= hist179 ( 31 downto 0 );
hist( 5791 downto 5760 ) <= hist180 ( 31 downto 0 );
hist( 5823 downto 5792 ) <= hist181 ( 31 downto 0 );
hist( 5855 downto 5824 ) <= hist182 ( 31 downto 0 );
hist( 5887 downto 5856 ) <= hist183 ( 31 downto 0 );
hist( 5919 downto 5888 ) <= hist184 ( 31 downto 0 );
hist( 5951 downto 5920 ) <= hist185 ( 31 downto 0 );
hist( 5983 downto 5952 ) <= hist186 ( 31 downto 0 );
hist( 6015 downto 5984 ) <= hist187 ( 31 downto 0 );
hist( 6047 downto 6016 ) <= hist188 ( 31 downto 0 );
hist( 6079 downto 6048 ) <= hist189 ( 31 downto 0 );
hist( 6111 downto 6080 ) <= hist190 ( 31 downto 0 );
hist( 6143 downto 6112 ) <= hist191 ( 31 downto 0 );
hist( 6175 downto 6144 ) <= hist192 ( 31 downto 0 );
hist( 6207 downto 6176 ) <= hist193 ( 31 downto 0 );
hist( 6239 downto 6208 ) <= hist194 ( 31 downto 0 );
hist( 6271 downto 6240 ) <= hist195 ( 31 downto 0 );
hist( 6303 downto 6272 ) <= hist196 ( 31 downto 0 );
hist( 6335 downto 6304 ) <= hist197 ( 31 downto 0 );
hist( 6367 downto 6336 ) <= hist198 ( 31 downto 0 );
hist( 6399 downto 6368 ) <= hist199 ( 31 downto 0 );
hist( 6431 downto 6400 ) <= hist200 ( 31 downto 0 );
hist( 6463 downto 6432 ) <= hist201 ( 31 downto 0 );
hist( 6495 downto 6464 ) <= hist202 ( 31 downto 0 );
hist( 6527 downto 6496 ) <= hist203 ( 31 downto 0 );
hist( 6559 downto 6528 ) <= hist204 ( 31 downto 0 );
hist( 6591 downto 6560 ) <= hist205 ( 31 downto 0 );
hist( 6623 downto 6592 ) <= hist206 ( 31 downto 0 );
hist( 6655 downto 6624 ) <= hist207 ( 31 downto 0 );
hist( 6687 downto 6656 ) <= hist208 ( 31 downto 0 );
hist( 6719 downto 6688 ) <= hist209 ( 31 downto 0 );
hist( 6751 downto 6720 ) <= hist210 ( 31 downto 0 );
hist( 6783 downto 6752 ) <= hist211 ( 31 downto 0 );
hist( 6815 downto 6784 ) <= hist212 ( 31 downto 0 );
hist( 6847 downto 6816 ) <= hist213 ( 31 downto 0 );
hist( 6879 downto 6848 ) <= hist214 ( 31 downto 0 );
hist( 6911 downto 6880 ) <= hist215 ( 31 downto 0 );
hist( 6943 downto 6912 ) <= hist216 ( 31 downto 0 );
hist( 6975 downto 6944 ) <= hist217 ( 31 downto 0 );
hist( 7007 downto 6976 ) <= hist218 ( 31 downto 0 );
hist( 7039 downto 7008 ) <= hist219 ( 31 downto 0 );
hist( 7071 downto 7040 ) <= hist220 ( 31 downto 0 );
hist( 7103 downto 7072 ) <= hist221 ( 31 downto 0 );
hist( 7135 downto 7104 ) <= hist222 ( 31 downto 0 );
hist( 7167 downto 7136 ) <= hist223 ( 31 downto 0 );
hist( 7199 downto 7168 ) <= hist224 ( 31 downto 0 );
hist( 7231 downto 7200 ) <= hist225 ( 31 downto 0 );
hist( 7263 downto 7232 ) <= hist226 ( 31 downto 0 );
hist( 7295 downto 7264 ) <= hist227 ( 31 downto 0 );
hist( 7327 downto 7296 ) <= hist228 ( 31 downto 0 );
hist( 7359 downto 7328 ) <= hist229 ( 31 downto 0 );
hist( 7391 downto 7360 ) <= hist230 ( 31 downto 0 );
hist( 7423 downto 7392 ) <= hist231 ( 31 downto 0 );
hist( 7455 downto 7424 ) <= hist232 ( 31 downto 0 );
hist( 7487 downto 7456 ) <= hist233 ( 31 downto 0 );
hist( 7519 downto 7488 ) <= hist234 ( 31 downto 0 );
hist( 7551 downto 7520 ) <= hist235 ( 31 downto 0 );
hist( 7583 downto 7552 ) <= hist236 ( 31 downto 0 );
hist( 7615 downto 7584 ) <= hist237 ( 31 downto 0 );
hist( 7647 downto 7616 ) <= hist238 ( 31 downto 0 );
hist( 7679 downto 7648 ) <= hist239 ( 31 downto 0 );
hist( 7711 downto 7680 ) <= hist240 ( 31 downto 0 );
hist( 7743 downto 7712 ) <= hist241 ( 31 downto 0 );
hist( 7775 downto 7744 ) <= hist242 ( 31 downto 0 );
hist( 7807 downto 7776 ) <= hist243 ( 31 downto 0 );
hist( 7839 downto 7808 ) <= hist244 ( 31 downto 0 );
hist( 7871 downto 7840 ) <= hist245 ( 31 downto 0 );
hist( 7903 downto 7872 ) <= hist246 ( 31 downto 0 );
hist( 7935 downto 7904 ) <= hist247 ( 31 downto 0 );
hist( 7967 downto 7936 ) <= hist248 ( 31 downto 0 );
hist( 7999 downto 7968 ) <= hist249 ( 31 downto 0 );
hist( 8031 downto 8000 ) <= hist250 ( 31 downto 0 );
hist( 8063 downto 8032 ) <= hist251 ( 31 downto 0 );
hist( 8095 downto 8064 ) <= hist252 ( 31 downto 0 );
hist( 8127 downto 8096 ) <= hist253 ( 31 downto 0 );
hist( 8159 downto 8128 ) <= hist254 ( 31 downto 0 );
hist( 8191 downto 8160 ) <= hist255 ( 31 downto 0 );
hist( 8223 downto 8192 ) <= hist256 ( 31 downto 0 );
hist( 8255 downto 8224 ) <= hist257 ( 31 downto 0 );
hist( 8287 downto 8256 ) <= hist258 ( 31 downto 0 );
hist( 8319 downto 8288 ) <= hist259 ( 31 downto 0 );
hist( 8351 downto 8320 ) <= hist260 ( 31 downto 0 );
hist( 8383 downto 8352 ) <= hist261 ( 31 downto 0 );
hist( 8415 downto 8384 ) <= hist262 ( 31 downto 0 );
hist( 8447 downto 8416 ) <= hist263 ( 31 downto 0 );
hist( 8479 downto 8448 ) <= hist264 ( 31 downto 0 );
hist( 8511 downto 8480 ) <= hist265 ( 31 downto 0 );
hist( 8543 downto 8512 ) <= hist266 ( 31 downto 0 );
hist( 8575 downto 8544 ) <= hist267 ( 31 downto 0 );
hist( 8607 downto 8576 ) <= hist268 ( 31 downto 0 );
hist( 8639 downto 8608 ) <= hist269 ( 31 downto 0 );
hist( 8671 downto 8640 ) <= hist270 ( 31 downto 0 );
hist( 8703 downto 8672 ) <= hist271 ( 31 downto 0 );
hist( 8735 downto 8704 ) <= hist272 ( 31 downto 0 );
hist( 8767 downto 8736 ) <= hist273 ( 31 downto 0 );
hist( 8799 downto 8768 ) <= hist274 ( 31 downto 0 );
hist( 8831 downto 8800 ) <= hist275 ( 31 downto 0 );
hist( 8863 downto 8832 ) <= hist276 ( 31 downto 0 );
hist( 8895 downto 8864 ) <= hist277 ( 31 downto 0 );
hist( 8927 downto 8896 ) <= hist278 ( 31 downto 0 );
hist( 8959 downto 8928 ) <= hist279 ( 31 downto 0 );
hist( 8991 downto 8960 ) <= hist280 ( 31 downto 0 );
hist( 9023 downto 8992 ) <= hist281 ( 31 downto 0 );
hist( 9055 downto 9024 ) <= hist282 ( 31 downto 0 );
hist( 9087 downto 9056 ) <= hist283 ( 31 downto 0 );
hist( 9119 downto 9088 ) <= hist284 ( 31 downto 0 );
hist( 9151 downto 9120 ) <= hist285 ( 31 downto 0 );
hist( 9183 downto 9152 ) <= hist286 ( 31 downto 0 );
hist( 9215 downto 9184 ) <= hist287 ( 31 downto 0 );
hist( 9247 downto 9216 ) <= hist288 ( 31 downto 0 );
hist( 9279 downto 9248 ) <= hist289 ( 31 downto 0 );
hist( 9311 downto 9280 ) <= hist290 ( 31 downto 0 );
hist( 9343 downto 9312 ) <= hist291 ( 31 downto 0 );
hist( 9375 downto 9344 ) <= hist292 ( 31 downto 0 );
hist( 9407 downto 9376 ) <= hist293 ( 31 downto 0 );
hist( 9439 downto 9408 ) <= hist294 ( 31 downto 0 );
hist( 9471 downto 9440 ) <= hist295 ( 31 downto 0 );
hist( 9503 downto 9472 ) <= hist296 ( 31 downto 0 );
hist( 9535 downto 9504 ) <= hist297 ( 31 downto 0 );
hist( 9567 downto 9536 ) <= hist298 ( 31 downto 0 );
hist( 9599 downto 9568 ) <= hist299 ( 31 downto 0 );
hist( 9631 downto 9600 ) <= hist300 ( 31 downto 0 );
hist( 9663 downto 9632 ) <= hist301 ( 31 downto 0 );
hist( 9695 downto 9664 ) <= hist302 ( 31 downto 0 );
hist( 9727 downto 9696 ) <= hist303 ( 31 downto 0 );
hist( 9759 downto 9728 ) <= hist304 ( 31 downto 0 );
hist( 9791 downto 9760 ) <= hist305 ( 31 downto 0 );
hist( 9823 downto 9792 ) <= hist306 ( 31 downto 0 );
hist( 9855 downto 9824 ) <= hist307 ( 31 downto 0 );
hist( 9887 downto 9856 ) <= hist308 ( 31 downto 0 );
hist( 9919 downto 9888 ) <= hist309 ( 31 downto 0 );
hist( 9951 downto 9920 ) <= hist310 ( 31 downto 0 );
hist( 9983 downto 9952 ) <= hist311 ( 31 downto 0 );
hist( 10015 downto 9984 ) <= hist312 ( 31 downto 0 );
hist( 10047 downto 10016 ) <= hist313 ( 31 downto 0 );
hist( 10079 downto 10048 ) <= hist314 ( 31 downto 0 );
hist( 10111 downto 10080 ) <= hist315 ( 31 downto 0 );
hist( 10143 downto 10112 ) <= hist316 ( 31 downto 0 );
hist( 10175 downto 10144 ) <= hist317 ( 31 downto 0 );
hist( 10207 downto 10176 ) <= hist318 ( 31 downto 0 );
hist( 10239 downto 10208 ) <= hist319 ( 31 downto 0 );
hist( 10271 downto 10240 ) <= hist320 ( 31 downto 0 );
hist( 10303 downto 10272 ) <= hist321 ( 31 downto 0 );
hist( 10335 downto 10304 ) <= hist322 ( 31 downto 0 );
hist( 10367 downto 10336 ) <= hist323 ( 31 downto 0 );
hist( 10399 downto 10368 ) <= hist324 ( 31 downto 0 );
hist( 10431 downto 10400 ) <= hist325 ( 31 downto 0 );
hist( 10463 downto 10432 ) <= hist326 ( 31 downto 0 );
hist( 10495 downto 10464 ) <= hist327 ( 31 downto 0 );
hist( 10527 downto 10496 ) <= hist328 ( 31 downto 0 );
hist( 10559 downto 10528 ) <= hist329 ( 31 downto 0 );
hist( 10591 downto 10560 ) <= hist330 ( 31 downto 0 );
hist( 10623 downto 10592 ) <= hist331 ( 31 downto 0 );
hist( 10655 downto 10624 ) <= hist332 ( 31 downto 0 );
hist( 10687 downto 10656 ) <= hist333 ( 31 downto 0 );
hist( 10719 downto 10688 ) <= hist334 ( 31 downto 0 );
hist( 10751 downto 10720 ) <= hist335 ( 31 downto 0 );
hist( 10783 downto 10752 ) <= hist336 ( 31 downto 0 );
hist( 10815 downto 10784 ) <= hist337 ( 31 downto 0 );
hist( 10847 downto 10816 ) <= hist338 ( 31 downto 0 );
hist( 10879 downto 10848 ) <= hist339 ( 31 downto 0 );
hist( 10911 downto 10880 ) <= hist340 ( 31 downto 0 );
hist( 10943 downto 10912 ) <= hist341 ( 31 downto 0 );
hist( 10975 downto 10944 ) <= hist342 ( 31 downto 0 );
hist( 11007 downto 10976 ) <= hist343 ( 31 downto 0 );
hist( 11039 downto 11008 ) <= hist344 ( 31 downto 0 );
hist( 11071 downto 11040 ) <= hist345 ( 31 downto 0 );
hist( 11103 downto 11072 ) <= hist346 ( 31 downto 0 );
hist( 11135 downto 11104 ) <= hist347 ( 31 downto 0 );
hist( 11167 downto 11136 ) <= hist348 ( 31 downto 0 );
hist( 11199 downto 11168 ) <= hist349 ( 31 downto 0 );
hist( 11231 downto 11200 ) <= hist350 ( 31 downto 0 );
hist( 11263 downto 11232 ) <= hist351 ( 31 downto 0 );
hist( 11295 downto 11264 ) <= hist352 ( 31 downto 0 );
hist( 11327 downto 11296 ) <= hist353 ( 31 downto 0 );
hist( 11359 downto 11328 ) <= hist354 ( 31 downto 0 );
hist( 11391 downto 11360 ) <= hist355 ( 31 downto 0 );
hist( 11423 downto 11392 ) <= hist356 ( 31 downto 0 );
hist( 11455 downto 11424 ) <= hist357 ( 31 downto 0 );
hist( 11487 downto 11456 ) <= hist358 ( 31 downto 0 );
hist( 11519 downto 11488 ) <= hist359 ( 31 downto 0 );
hist( 11551 downto 11520 ) <= hist360 ( 31 downto 0 );
hist( 11583 downto 11552 ) <= hist361 ( 31 downto 0 );
hist( 11615 downto 11584 ) <= hist362 ( 31 downto 0 );
hist( 11647 downto 11616 ) <= hist363 ( 31 downto 0 );
hist( 11679 downto 11648 ) <= hist364 ( 31 downto 0 );
hist( 11711 downto 11680 ) <= hist365 ( 31 downto 0 );
hist( 11743 downto 11712 ) <= hist366 ( 31 downto 0 );
hist( 11775 downto 11744 ) <= hist367 ( 31 downto 0 );
hist( 11807 downto 11776 ) <= hist368 ( 31 downto 0 );
hist( 11839 downto 11808 ) <= hist369 ( 31 downto 0 );
hist( 11871 downto 11840 ) <= hist370 ( 31 downto 0 );
hist( 11903 downto 11872 ) <= hist371 ( 31 downto 0 );
hist( 11935 downto 11904 ) <= hist372 ( 31 downto 0 );
hist( 11967 downto 11936 ) <= hist373 ( 31 downto 0 );
hist( 11999 downto 11968 ) <= hist374 ( 31 downto 0 );
hist( 12031 downto 12000 ) <= hist375 ( 31 downto 0 );
hist( 12063 downto 12032 ) <= hist376 ( 31 downto 0 );
hist( 12095 downto 12064 ) <= hist377 ( 31 downto 0 );
hist( 12127 downto 12096 ) <= hist378 ( 31 downto 0 );
hist( 12159 downto 12128 ) <= hist379 ( 31 downto 0 );
hist( 12191 downto 12160 ) <= hist380 ( 31 downto 0 );
hist( 12223 downto 12192 ) <= hist381 ( 31 downto 0 );
hist( 12255 downto 12224 ) <= hist382 ( 31 downto 0 );
hist( 12287 downto 12256 ) <= hist383 ( 31 downto 0 );
hist( 12319 downto 12288 ) <= hist384 ( 31 downto 0 );
hist( 12351 downto 12320 ) <= hist385 ( 31 downto 0 );
hist( 12383 downto 12352 ) <= hist386 ( 31 downto 0 );
hist( 12415 downto 12384 ) <= hist387 ( 31 downto 0 );
hist( 12447 downto 12416 ) <= hist388 ( 31 downto 0 );
hist( 12479 downto 12448 ) <= hist389 ( 31 downto 0 );
hist( 12511 downto 12480 ) <= hist390 ( 31 downto 0 );
hist( 12543 downto 12512 ) <= hist391 ( 31 downto 0 );
hist( 12575 downto 12544 ) <= hist392 ( 31 downto 0 );
hist( 12607 downto 12576 ) <= hist393 ( 31 downto 0 );
hist( 12639 downto 12608 ) <= hist394 ( 31 downto 0 );
hist( 12671 downto 12640 ) <= hist395 ( 31 downto 0 );
hist( 12703 downto 12672 ) <= hist396 ( 31 downto 0 );
hist( 12735 downto 12704 ) <= hist397 ( 31 downto 0 );
hist( 12767 downto 12736 ) <= hist398 ( 31 downto 0 );
hist( 12799 downto 12768 ) <= hist399 ( 31 downto 0 );
hist( 12831 downto 12800 ) <= hist400 ( 31 downto 0 );
hist( 12863 downto 12832 ) <= hist401 ( 31 downto 0 );
hist( 12895 downto 12864 ) <= hist402 ( 31 downto 0 );
hist( 12927 downto 12896 ) <= hist403 ( 31 downto 0 );
hist( 12959 downto 12928 ) <= hist404 ( 31 downto 0 );
hist( 12991 downto 12960 ) <= hist405 ( 31 downto 0 );
hist( 13023 downto 12992 ) <= hist406 ( 31 downto 0 );
hist( 13055 downto 13024 ) <= hist407 ( 31 downto 0 );
hist( 13087 downto 13056 ) <= hist408 ( 31 downto 0 );
hist( 13119 downto 13088 ) <= hist409 ( 31 downto 0 );
hist( 13151 downto 13120 ) <= hist410 ( 31 downto 0 );
hist( 13183 downto 13152 ) <= hist411 ( 31 downto 0 );
hist( 13215 downto 13184 ) <= hist412 ( 31 downto 0 );
hist( 13247 downto 13216 ) <= hist413 ( 31 downto 0 );
hist( 13279 downto 13248 ) <= hist414 ( 31 downto 0 );
hist( 13311 downto 13280 ) <= hist415 ( 31 downto 0 );
hist( 13343 downto 13312 ) <= hist416 ( 31 downto 0 );
hist( 13375 downto 13344 ) <= hist417 ( 31 downto 0 );
hist( 13407 downto 13376 ) <= hist418 ( 31 downto 0 );
hist( 13439 downto 13408 ) <= hist419 ( 31 downto 0 );
hist( 13471 downto 13440 ) <= hist420 ( 31 downto 0 );
hist( 13503 downto 13472 ) <= hist421 ( 31 downto 0 );
hist( 13535 downto 13504 ) <= hist422 ( 31 downto 0 );
hist( 13567 downto 13536 ) <= hist423 ( 31 downto 0 );
hist( 13599 downto 13568 ) <= hist424 ( 31 downto 0 );
hist( 13631 downto 13600 ) <= hist425 ( 31 downto 0 );
hist( 13663 downto 13632 ) <= hist426 ( 31 downto 0 );
hist( 13695 downto 13664 ) <= hist427 ( 31 downto 0 );
hist( 13727 downto 13696 ) <= hist428 ( 31 downto 0 );
hist( 13759 downto 13728 ) <= hist429 ( 31 downto 0 );
hist( 13791 downto 13760 ) <= hist430 ( 31 downto 0 );
hist( 13823 downto 13792 ) <= hist431 ( 31 downto 0 );
hist( 13855 downto 13824 ) <= hist432 ( 31 downto 0 );
hist( 13887 downto 13856 ) <= hist433 ( 31 downto 0 );
hist( 13919 downto 13888 ) <= hist434 ( 31 downto 0 );
hist( 13951 downto 13920 ) <= hist435 ( 31 downto 0 );
hist( 13983 downto 13952 ) <= hist436 ( 31 downto 0 );
hist( 14015 downto 13984 ) <= hist437 ( 31 downto 0 );
hist( 14047 downto 14016 ) <= hist438 ( 31 downto 0 );
hist( 14079 downto 14048 ) <= hist439 ( 31 downto 0 );
hist( 14111 downto 14080 ) <= hist440 ( 31 downto 0 );
hist( 14143 downto 14112 ) <= hist441 ( 31 downto 0 );
hist( 14175 downto 14144 ) <= hist442 ( 31 downto 0 );
hist( 14207 downto 14176 ) <= hist443 ( 31 downto 0 );
hist( 14239 downto 14208 ) <= hist444 ( 31 downto 0 );
hist( 14271 downto 14240 ) <= hist445 ( 31 downto 0 );
hist( 14303 downto 14272 ) <= hist446 ( 31 downto 0 );
hist( 14335 downto 14304 ) <= hist447 ( 31 downto 0 );
hist( 14367 downto 14336 ) <= hist448 ( 31 downto 0 );
hist( 14399 downto 14368 ) <= hist449 ( 31 downto 0 );
hist( 14431 downto 14400 ) <= hist450 ( 31 downto 0 );
hist( 14463 downto 14432 ) <= hist451 ( 31 downto 0 );
hist( 14495 downto 14464 ) <= hist452 ( 31 downto 0 );
hist( 14527 downto 14496 ) <= hist453 ( 31 downto 0 );
hist( 14559 downto 14528 ) <= hist454 ( 31 downto 0 );
hist( 14591 downto 14560 ) <= hist455 ( 31 downto 0 );
hist( 14623 downto 14592 ) <= hist456 ( 31 downto 0 );
hist( 14655 downto 14624 ) <= hist457 ( 31 downto 0 );
hist( 14687 downto 14656 ) <= hist458 ( 31 downto 0 );
hist( 14719 downto 14688 ) <= hist459 ( 31 downto 0 );
hist( 14751 downto 14720 ) <= hist460 ( 31 downto 0 );
hist( 14783 downto 14752 ) <= hist461 ( 31 downto 0 );
hist( 14815 downto 14784 ) <= hist462 ( 31 downto 0 );
hist( 14847 downto 14816 ) <= hist463 ( 31 downto 0 );
hist( 14879 downto 14848 ) <= hist464 ( 31 downto 0 );
hist( 14911 downto 14880 ) <= hist465 ( 31 downto 0 );
hist( 14943 downto 14912 ) <= hist466 ( 31 downto 0 );
hist( 14975 downto 14944 ) <= hist467 ( 31 downto 0 );
hist( 15007 downto 14976 ) <= hist468 ( 31 downto 0 );
hist( 15039 downto 15008 ) <= hist469 ( 31 downto 0 );
hist( 15071 downto 15040 ) <= hist470 ( 31 downto 0 );
hist( 15103 downto 15072 ) <= hist471 ( 31 downto 0 );
hist( 15135 downto 15104 ) <= hist472 ( 31 downto 0 );
hist( 15167 downto 15136 ) <= hist473 ( 31 downto 0 );
hist( 15199 downto 15168 ) <= hist474 ( 31 downto 0 );
hist( 15231 downto 15200 ) <= hist475 ( 31 downto 0 );
hist( 15263 downto 15232 ) <= hist476 ( 31 downto 0 );
hist( 15295 downto 15264 ) <= hist477 ( 31 downto 0 );
hist( 15327 downto 15296 ) <= hist478 ( 31 downto 0 );
hist( 15359 downto 15328 ) <= hist479 ( 31 downto 0 );
hist( 15391 downto 15360 ) <= hist480 ( 31 downto 0 );
hist( 15423 downto 15392 ) <= hist481 ( 31 downto 0 );
hist( 15455 downto 15424 ) <= hist482 ( 31 downto 0 );
hist( 15487 downto 15456 ) <= hist483 ( 31 downto 0 );
hist( 15519 downto 15488 ) <= hist484 ( 31 downto 0 );
hist( 15551 downto 15520 ) <= hist485 ( 31 downto 0 );
hist( 15583 downto 15552 ) <= hist486 ( 31 downto 0 );
hist( 15615 downto 15584 ) <= hist487 ( 31 downto 0 );
hist( 15647 downto 15616 ) <= hist488 ( 31 downto 0 );
hist( 15679 downto 15648 ) <= hist489 ( 31 downto 0 );
hist( 15711 downto 15680 ) <= hist490 ( 31 downto 0 );
hist( 15743 downto 15712 ) <= hist491 ( 31 downto 0 );
hist( 15775 downto 15744 ) <= hist492 ( 31 downto 0 );
hist( 15807 downto 15776 ) <= hist493 ( 31 downto 0 );
hist( 15839 downto 15808 ) <= hist494 ( 31 downto 0 );
hist( 15871 downto 15840 ) <= hist495 ( 31 downto 0 );
hist( 15903 downto 15872 ) <= hist496 ( 31 downto 0 );
hist( 15935 downto 15904 ) <= hist497 ( 31 downto 0 );
hist( 15967 downto 15936 ) <= hist498 ( 31 downto 0 );
hist( 15999 downto 15968 ) <= hist499 ( 31 downto 0 );
hist( 16031 downto 16000 ) <= hist500 ( 31 downto 0 );
hist( 16063 downto 16032 ) <= hist501 ( 31 downto 0 );
hist( 16095 downto 16064 ) <= hist502 ( 31 downto 0 );
hist( 16127 downto 16096 ) <= hist503 ( 31 downto 0 );
hist( 16159 downto 16128 ) <= hist504 ( 31 downto 0 );
hist( 16191 downto 16160 ) <= hist505 ( 31 downto 0 );
hist( 16223 downto 16192 ) <= hist506 ( 31 downto 0 );
hist( 16255 downto 16224 ) <= hist507 ( 31 downto 0 );
hist( 16287 downto 16256 ) <= hist508 ( 31 downto 0 );
hist( 16319 downto 16288 ) <= hist509 ( 31 downto 0 );
hist( 16351 downto 16320 ) <= hist510 ( 31 downto 0 );
hist( 16383 downto 16352 ) <= hist511 ( 31 downto 0 );
hist( 16415 downto 16384 ) <= hist512 ( 31 downto 0 );
hist( 16447 downto 16416 ) <= hist513 ( 31 downto 0 );
hist( 16479 downto 16448 ) <= hist514 ( 31 downto 0 );
hist( 16511 downto 16480 ) <= hist515 ( 31 downto 0 );
hist( 16543 downto 16512 ) <= hist516 ( 31 downto 0 );
hist( 16575 downto 16544 ) <= hist517 ( 31 downto 0 );
hist( 16607 downto 16576 ) <= hist518 ( 31 downto 0 );
hist( 16639 downto 16608 ) <= hist519 ( 31 downto 0 );
hist( 16671 downto 16640 ) <= hist520 ( 31 downto 0 );
hist( 16703 downto 16672 ) <= hist521 ( 31 downto 0 );
hist( 16735 downto 16704 ) <= hist522 ( 31 downto 0 );
hist( 16767 downto 16736 ) <= hist523 ( 31 downto 0 );
hist( 16799 downto 16768 ) <= hist524 ( 31 downto 0 );
hist( 16831 downto 16800 ) <= hist525 ( 31 downto 0 );
hist( 16863 downto 16832 ) <= hist526 ( 31 downto 0 );
hist( 16895 downto 16864 ) <= hist527 ( 31 downto 0 );
hist( 16927 downto 16896 ) <= hist528 ( 31 downto 0 );
hist( 16959 downto 16928 ) <= hist529 ( 31 downto 0 );
hist( 16991 downto 16960 ) <= hist530 ( 31 downto 0 );
hist( 17023 downto 16992 ) <= hist531 ( 31 downto 0 );
hist( 17055 downto 17024 ) <= hist532 ( 31 downto 0 );
hist( 17087 downto 17056 ) <= hist533 ( 31 downto 0 );
hist( 17119 downto 17088 ) <= hist534 ( 31 downto 0 );
hist( 17151 downto 17120 ) <= hist535 ( 31 downto 0 );
hist( 17183 downto 17152 ) <= hist536 ( 31 downto 0 );
hist( 17215 downto 17184 ) <= hist537 ( 31 downto 0 );
hist( 17247 downto 17216 ) <= hist538 ( 31 downto 0 );
hist( 17279 downto 17248 ) <= hist539 ( 31 downto 0 );
hist( 17311 downto 17280 ) <= hist540 ( 31 downto 0 );
hist( 17343 downto 17312 ) <= hist541 ( 31 downto 0 );
hist( 17375 downto 17344 ) <= hist542 ( 31 downto 0 );
hist( 17407 downto 17376 ) <= hist543 ( 31 downto 0 );
hist( 17439 downto 17408 ) <= hist544 ( 31 downto 0 );
hist( 17471 downto 17440 ) <= hist545 ( 31 downto 0 );
hist( 17503 downto 17472 ) <= hist546 ( 31 downto 0 );
hist( 17535 downto 17504 ) <= hist547 ( 31 downto 0 );
hist( 17567 downto 17536 ) <= hist548 ( 31 downto 0 );
hist( 17599 downto 17568 ) <= hist549 ( 31 downto 0 );
hist( 17631 downto 17600 ) <= hist550 ( 31 downto 0 );
hist( 17663 downto 17632 ) <= hist551 ( 31 downto 0 );
hist( 17695 downto 17664 ) <= hist552 ( 31 downto 0 );
hist( 17727 downto 17696 ) <= hist553 ( 31 downto 0 );
hist( 17759 downto 17728 ) <= hist554 ( 31 downto 0 );
hist( 17791 downto 17760 ) <= hist555 ( 31 downto 0 );
hist( 17823 downto 17792 ) <= hist556 ( 31 downto 0 );
hist( 17855 downto 17824 ) <= hist557 ( 31 downto 0 );
hist( 17887 downto 17856 ) <= hist558 ( 31 downto 0 );
hist( 17919 downto 17888 ) <= hist559 ( 31 downto 0 );
hist( 17951 downto 17920 ) <= hist560 ( 31 downto 0 );
hist( 17983 downto 17952 ) <= hist561 ( 31 downto 0 );
hist( 18015 downto 17984 ) <= hist562 ( 31 downto 0 );
hist( 18047 downto 18016 ) <= hist563 ( 31 downto 0 );
hist( 18079 downto 18048 ) <= hist564 ( 31 downto 0 );
hist( 18111 downto 18080 ) <= hist565 ( 31 downto 0 );
hist( 18143 downto 18112 ) <= hist566 ( 31 downto 0 );
hist( 18175 downto 18144 ) <= hist567 ( 31 downto 0 );
hist( 18207 downto 18176 ) <= hist568 ( 31 downto 0 );
hist( 18239 downto 18208 ) <= hist569 ( 31 downto 0 );
hist( 18271 downto 18240 ) <= hist570 ( 31 downto 0 );
hist( 18303 downto 18272 ) <= hist571 ( 31 downto 0 );
hist( 18335 downto 18304 ) <= hist572 ( 31 downto 0 );
hist( 18367 downto 18336 ) <= hist573 ( 31 downto 0 );
hist( 18399 downto 18368 ) <= hist574 ( 31 downto 0 );
hist( 18431 downto 18400 ) <= hist575 ( 31 downto 0 );
hist( 18463 downto 18432 ) <= hist576 ( 31 downto 0 );
hist( 18495 downto 18464 ) <= hist577 ( 31 downto 0 );
hist( 18527 downto 18496 ) <= hist578 ( 31 downto 0 );
hist( 18559 downto 18528 ) <= hist579 ( 31 downto 0 );
hist( 18591 downto 18560 ) <= hist580 ( 31 downto 0 );
hist( 18623 downto 18592 ) <= hist581 ( 31 downto 0 );
hist( 18655 downto 18624 ) <= hist582 ( 31 downto 0 );
hist( 18687 downto 18656 ) <= hist583 ( 31 downto 0 );
hist( 18719 downto 18688 ) <= hist584 ( 31 downto 0 );
hist( 18751 downto 18720 ) <= hist585 ( 31 downto 0 );
hist( 18783 downto 18752 ) <= hist586 ( 31 downto 0 );
hist( 18815 downto 18784 ) <= hist587 ( 31 downto 0 );
hist( 18847 downto 18816 ) <= hist588 ( 31 downto 0 );
hist( 18879 downto 18848 ) <= hist589 ( 31 downto 0 );
hist( 18911 downto 18880 ) <= hist590 ( 31 downto 0 );
hist( 18943 downto 18912 ) <= hist591 ( 31 downto 0 );
hist( 18975 downto 18944 ) <= hist592 ( 31 downto 0 );
hist( 19007 downto 18976 ) <= hist593 ( 31 downto 0 );
hist( 19039 downto 19008 ) <= hist594 ( 31 downto 0 );
hist( 19071 downto 19040 ) <= hist595 ( 31 downto 0 );
hist( 19103 downto 19072 ) <= hist596 ( 31 downto 0 );
hist( 19135 downto 19104 ) <= hist597 ( 31 downto 0 );
hist( 19167 downto 19136 ) <= hist598 ( 31 downto 0 );
hist( 19199 downto 19168 ) <= hist599 ( 31 downto 0 );
hist( 19231 downto 19200 ) <= hist600 ( 31 downto 0 );
hist( 19263 downto 19232 ) <= hist601 ( 31 downto 0 );
hist( 19295 downto 19264 ) <= hist602 ( 31 downto 0 );
hist( 19327 downto 19296 ) <= hist603 ( 31 downto 0 );
hist( 19359 downto 19328 ) <= hist604 ( 31 downto 0 );
hist( 19391 downto 19360 ) <= hist605 ( 31 downto 0 );
hist( 19423 downto 19392 ) <= hist606 ( 31 downto 0 );
hist( 19455 downto 19424 ) <= hist607 ( 31 downto 0 );
hist( 19487 downto 19456 ) <= hist608 ( 31 downto 0 );
hist( 19519 downto 19488 ) <= hist609 ( 31 downto 0 );
hist( 19551 downto 19520 ) <= hist610 ( 31 downto 0 );
hist( 19583 downto 19552 ) <= hist611 ( 31 downto 0 );
hist( 19615 downto 19584 ) <= hist612 ( 31 downto 0 );
hist( 19647 downto 19616 ) <= hist613 ( 31 downto 0 );
hist( 19679 downto 19648 ) <= hist614 ( 31 downto 0 );
hist( 19711 downto 19680 ) <= hist615 ( 31 downto 0 );
hist( 19743 downto 19712 ) <= hist616 ( 31 downto 0 );
hist( 19775 downto 19744 ) <= hist617 ( 31 downto 0 );
hist( 19807 downto 19776 ) <= hist618 ( 31 downto 0 );
hist( 19839 downto 19808 ) <= hist619 ( 31 downto 0 );
hist( 19871 downto 19840 ) <= hist620 ( 31 downto 0 );
hist( 19903 downto 19872 ) <= hist621 ( 31 downto 0 );
hist( 19935 downto 19904 ) <= hist622 ( 31 downto 0 );
hist( 19967 downto 19936 ) <= hist623 ( 31 downto 0 );
hist( 19999 downto 19968 ) <= hist624 ( 31 downto 0 );
hist( 20031 downto 20000 ) <= hist625 ( 31 downto 0 );
hist( 20063 downto 20032 ) <= hist626 ( 31 downto 0 );
hist( 20095 downto 20064 ) <= hist627 ( 31 downto 0 );
hist( 20127 downto 20096 ) <= hist628 ( 31 downto 0 );
hist( 20159 downto 20128 ) <= hist629 ( 31 downto 0 );
hist( 20191 downto 20160 ) <= hist630 ( 31 downto 0 );
hist( 20223 downto 20192 ) <= hist631 ( 31 downto 0 );
hist( 20255 downto 20224 ) <= hist632 ( 31 downto 0 );
hist( 20287 downto 20256 ) <= hist633 ( 31 downto 0 );
hist( 20319 downto 20288 ) <= hist634 ( 31 downto 0 );
hist( 20351 downto 20320 ) <= hist635 ( 31 downto 0 );
hist( 20383 downto 20352 ) <= hist636 ( 31 downto 0 );
hist( 20415 downto 20384 ) <= hist637 ( 31 downto 0 );
hist( 20447 downto 20416 ) <= hist638 ( 31 downto 0 );
hist( 20479 downto 20448 ) <= hist639 ( 31 downto 0 );
hist( 20511 downto 20480 ) <= hist640 ( 31 downto 0 );
hist( 20543 downto 20512 ) <= hist641 ( 31 downto 0 );
hist( 20575 downto 20544 ) <= hist642 ( 31 downto 0 );
hist( 20607 downto 20576 ) <= hist643 ( 31 downto 0 );
hist( 20639 downto 20608 ) <= hist644 ( 31 downto 0 );
hist( 20671 downto 20640 ) <= hist645 ( 31 downto 0 );
hist( 20703 downto 20672 ) <= hist646 ( 31 downto 0 );
hist( 20735 downto 20704 ) <= hist647 ( 31 downto 0 );
hist( 20767 downto 20736 ) <= hist648 ( 31 downto 0 );
hist( 20799 downto 20768 ) <= hist649 ( 31 downto 0 );
hist( 20831 downto 20800 ) <= hist650 ( 31 downto 0 );
hist( 20863 downto 20832 ) <= hist651 ( 31 downto 0 );
hist( 20895 downto 20864 ) <= hist652 ( 31 downto 0 );
hist( 20927 downto 20896 ) <= hist653 ( 31 downto 0 );
hist( 20959 downto 20928 ) <= hist654 ( 31 downto 0 );
hist( 20991 downto 20960 ) <= hist655 ( 31 downto 0 );
hist( 21023 downto 20992 ) <= hist656 ( 31 downto 0 );
hist( 21055 downto 21024 ) <= hist657 ( 31 downto 0 );
hist( 21087 downto 21056 ) <= hist658 ( 31 downto 0 );
hist( 21119 downto 21088 ) <= hist659 ( 31 downto 0 );
hist( 21151 downto 21120 ) <= hist660 ( 31 downto 0 );
hist( 21183 downto 21152 ) <= hist661 ( 31 downto 0 );
hist( 21215 downto 21184 ) <= hist662 ( 31 downto 0 );
hist( 21247 downto 21216 ) <= hist663 ( 31 downto 0 );
hist( 21279 downto 21248 ) <= hist664 ( 31 downto 0 );
hist( 21311 downto 21280 ) <= hist665 ( 31 downto 0 );
hist( 21343 downto 21312 ) <= hist666 ( 31 downto 0 );
hist( 21375 downto 21344 ) <= hist667 ( 31 downto 0 );
hist( 21407 downto 21376 ) <= hist668 ( 31 downto 0 );
hist( 21439 downto 21408 ) <= hist669 ( 31 downto 0 );
hist( 21471 downto 21440 ) <= hist670 ( 31 downto 0 );
hist( 21503 downto 21472 ) <= hist671 ( 31 downto 0 );
hist( 21535 downto 21504 ) <= hist672 ( 31 downto 0 );
hist( 21567 downto 21536 ) <= hist673 ( 31 downto 0 );
hist( 21599 downto 21568 ) <= hist674 ( 31 downto 0 );
hist( 21631 downto 21600 ) <= hist675 ( 31 downto 0 );
hist( 21663 downto 21632 ) <= hist676 ( 31 downto 0 );
hist( 21695 downto 21664 ) <= hist677 ( 31 downto 0 );
hist( 21727 downto 21696 ) <= hist678 ( 31 downto 0 );
hist( 21759 downto 21728 ) <= hist679 ( 31 downto 0 );
hist( 21791 downto 21760 ) <= hist680 ( 31 downto 0 );
hist( 21823 downto 21792 ) <= hist681 ( 31 downto 0 );
hist( 21855 downto 21824 ) <= hist682 ( 31 downto 0 );
hist( 21887 downto 21856 ) <= hist683 ( 31 downto 0 );
hist( 21919 downto 21888 ) <= hist684 ( 31 downto 0 );
hist( 21951 downto 21920 ) <= hist685 ( 31 downto 0 );
hist( 21983 downto 21952 ) <= hist686 ( 31 downto 0 );
hist( 22015 downto 21984 ) <= hist687 ( 31 downto 0 );
hist( 22047 downto 22016 ) <= hist688 ( 31 downto 0 );
hist( 22079 downto 22048 ) <= hist689 ( 31 downto 0 );
hist( 22111 downto 22080 ) <= hist690 ( 31 downto 0 );
hist( 22143 downto 22112 ) <= hist691 ( 31 downto 0 );
hist( 22175 downto 22144 ) <= hist692 ( 31 downto 0 );
hist( 22207 downto 22176 ) <= hist693 ( 31 downto 0 );
hist( 22239 downto 22208 ) <= hist694 ( 31 downto 0 );
hist( 22271 downto 22240 ) <= hist695 ( 31 downto 0 );
hist( 22303 downto 22272 ) <= hist696 ( 31 downto 0 );
hist( 22335 downto 22304 ) <= hist697 ( 31 downto 0 );
hist( 22367 downto 22336 ) <= hist698 ( 31 downto 0 );
hist( 22399 downto 22368 ) <= hist699 ( 31 downto 0 );
hist( 22431 downto 22400 ) <= hist700 ( 31 downto 0 );
hist( 22463 downto 22432 ) <= hist701 ( 31 downto 0 );
hist( 22495 downto 22464 ) <= hist702 ( 31 downto 0 );
hist( 22527 downto 22496 ) <= hist703 ( 31 downto 0 );
hist( 22559 downto 22528 ) <= hist704 ( 31 downto 0 );
hist( 22591 downto 22560 ) <= hist705 ( 31 downto 0 );
hist( 22623 downto 22592 ) <= hist706 ( 31 downto 0 );
hist( 22655 downto 22624 ) <= hist707 ( 31 downto 0 );
hist( 22687 downto 22656 ) <= hist708 ( 31 downto 0 );
hist( 22719 downto 22688 ) <= hist709 ( 31 downto 0 );
hist( 22751 downto 22720 ) <= hist710 ( 31 downto 0 );
hist( 22783 downto 22752 ) <= hist711 ( 31 downto 0 );
hist( 22815 downto 22784 ) <= hist712 ( 31 downto 0 );
hist( 22847 downto 22816 ) <= hist713 ( 31 downto 0 );
hist( 22879 downto 22848 ) <= hist714 ( 31 downto 0 );
hist( 22911 downto 22880 ) <= hist715 ( 31 downto 0 );
hist( 22943 downto 22912 ) <= hist716 ( 31 downto 0 );
hist( 22975 downto 22944 ) <= hist717 ( 31 downto 0 );
hist( 23007 downto 22976 ) <= hist718 ( 31 downto 0 );
hist( 23039 downto 23008 ) <= hist719 ( 31 downto 0 );
hist( 23071 downto 23040 ) <= hist720 ( 31 downto 0 );
hist( 23103 downto 23072 ) <= hist721 ( 31 downto 0 );
hist( 23135 downto 23104 ) <= hist722 ( 31 downto 0 );
hist( 23167 downto 23136 ) <= hist723 ( 31 downto 0 );
hist( 23199 downto 23168 ) <= hist724 ( 31 downto 0 );
hist( 23231 downto 23200 ) <= hist725 ( 31 downto 0 );
hist( 23263 downto 23232 ) <= hist726 ( 31 downto 0 );
hist( 23295 downto 23264 ) <= hist727 ( 31 downto 0 );
hist( 23327 downto 23296 ) <= hist728 ( 31 downto 0 );
hist( 23359 downto 23328 ) <= hist729 ( 31 downto 0 );
hist( 23391 downto 23360 ) <= hist730 ( 31 downto 0 );
hist( 23423 downto 23392 ) <= hist731 ( 31 downto 0 );
hist( 23455 downto 23424 ) <= hist732 ( 31 downto 0 );
hist( 23487 downto 23456 ) <= hist733 ( 31 downto 0 );
hist( 23519 downto 23488 ) <= hist734 ( 31 downto 0 );
hist( 23551 downto 23520 ) <= hist735 ( 31 downto 0 );
hist( 23583 downto 23552 ) <= hist736 ( 31 downto 0 );
hist( 23615 downto 23584 ) <= hist737 ( 31 downto 0 );
hist( 23647 downto 23616 ) <= hist738 ( 31 downto 0 );
hist( 23679 downto 23648 ) <= hist739 ( 31 downto 0 );
hist( 23711 downto 23680 ) <= hist740 ( 31 downto 0 );
hist( 23743 downto 23712 ) <= hist741 ( 31 downto 0 );
hist( 23775 downto 23744 ) <= hist742 ( 31 downto 0 );
hist( 23807 downto 23776 ) <= hist743 ( 31 downto 0 );
hist( 23839 downto 23808 ) <= hist744 ( 31 downto 0 );
hist( 23871 downto 23840 ) <= hist745 ( 31 downto 0 );
hist( 23903 downto 23872 ) <= hist746 ( 31 downto 0 );
hist( 23935 downto 23904 ) <= hist747 ( 31 downto 0 );
hist( 23967 downto 23936 ) <= hist748 ( 31 downto 0 );
hist( 23999 downto 23968 ) <= hist749 ( 31 downto 0 );
hist( 24031 downto 24000 ) <= hist750 ( 31 downto 0 );
hist( 24063 downto 24032 ) <= hist751 ( 31 downto 0 );
hist( 24095 downto 24064 ) <= hist752 ( 31 downto 0 );
hist( 24127 downto 24096 ) <= hist753 ( 31 downto 0 );
hist( 24159 downto 24128 ) <= hist754 ( 31 downto 0 );
hist( 24191 downto 24160 ) <= hist755 ( 31 downto 0 );
hist( 24223 downto 24192 ) <= hist756 ( 31 downto 0 );
hist( 24255 downto 24224 ) <= hist757 ( 31 downto 0 );
hist( 24287 downto 24256 ) <= hist758 ( 31 downto 0 );
hist( 24319 downto 24288 ) <= hist759 ( 31 downto 0 );
hist( 24351 downto 24320 ) <= hist760 ( 31 downto 0 );
hist( 24383 downto 24352 ) <= hist761 ( 31 downto 0 );
hist( 24415 downto 24384 ) <= hist762 ( 31 downto 0 );
hist( 24447 downto 24416 ) <= hist763 ( 31 downto 0 );
hist( 24479 downto 24448 ) <= hist764 ( 31 downto 0 );
hist( 24511 downto 24480 ) <= hist765 ( 31 downto 0 );
hist( 24543 downto 24512 ) <= hist766 ( 31 downto 0 );
hist( 24575 downto 24544 ) <= hist767 ( 31 downto 0 );
hist( 24607 downto 24576 ) <= hist768 ( 31 downto 0 );
hist( 24639 downto 24608 ) <= hist769 ( 31 downto 0 );
hist( 24671 downto 24640 ) <= hist770 ( 31 downto 0 );
hist( 24703 downto 24672 ) <= hist771 ( 31 downto 0 );
hist( 24735 downto 24704 ) <= hist772 ( 31 downto 0 );
hist( 24767 downto 24736 ) <= hist773 ( 31 downto 0 );
hist( 24799 downto 24768 ) <= hist774 ( 31 downto 0 );
hist( 24831 downto 24800 ) <= hist775 ( 31 downto 0 );
hist( 24863 downto 24832 ) <= hist776 ( 31 downto 0 );
hist( 24895 downto 24864 ) <= hist777 ( 31 downto 0 );
hist( 24927 downto 24896 ) <= hist778 ( 31 downto 0 );
hist( 24959 downto 24928 ) <= hist779 ( 31 downto 0 );
hist( 24991 downto 24960 ) <= hist780 ( 31 downto 0 );
hist( 25023 downto 24992 ) <= hist781 ( 31 downto 0 );
hist( 25055 downto 25024 ) <= hist782 ( 31 downto 0 );
hist( 25087 downto 25056 ) <= hist783 ( 31 downto 0 );
hist( 25119 downto 25088 ) <= hist784 ( 31 downto 0 );
hist( 25151 downto 25120 ) <= hist785 ( 31 downto 0 );
hist( 25183 downto 25152 ) <= hist786 ( 31 downto 0 );
hist( 25215 downto 25184 ) <= hist787 ( 31 downto 0 );
hist( 25247 downto 25216 ) <= hist788 ( 31 downto 0 );
hist( 25279 downto 25248 ) <= hist789 ( 31 downto 0 );
hist( 25311 downto 25280 ) <= hist790 ( 31 downto 0 );
hist( 25343 downto 25312 ) <= hist791 ( 31 downto 0 );
hist( 25375 downto 25344 ) <= hist792 ( 31 downto 0 );
hist( 25407 downto 25376 ) <= hist793 ( 31 downto 0 );
hist( 25439 downto 25408 ) <= hist794 ( 31 downto 0 );
hist( 25471 downto 25440 ) <= hist795 ( 31 downto 0 );
hist( 25503 downto 25472 ) <= hist796 ( 31 downto 0 );
hist( 25535 downto 25504 ) <= hist797 ( 31 downto 0 );
hist( 25567 downto 25536 ) <= hist798 ( 31 downto 0 );
hist( 25599 downto 25568 ) <= hist799 ( 31 downto 0 );
hist( 25631 downto 25600 ) <= hist800 ( 31 downto 0 );
hist( 25663 downto 25632 ) <= hist801 ( 31 downto 0 );
hist( 25695 downto 25664 ) <= hist802 ( 31 downto 0 );
hist( 25727 downto 25696 ) <= hist803 ( 31 downto 0 );
hist( 25759 downto 25728 ) <= hist804 ( 31 downto 0 );
hist( 25791 downto 25760 ) <= hist805 ( 31 downto 0 );
hist( 25823 downto 25792 ) <= hist806 ( 31 downto 0 );
hist( 25855 downto 25824 ) <= hist807 ( 31 downto 0 );
hist( 25887 downto 25856 ) <= hist808 ( 31 downto 0 );
hist( 25919 downto 25888 ) <= hist809 ( 31 downto 0 );
hist( 25951 downto 25920 ) <= hist810 ( 31 downto 0 );
hist( 25983 downto 25952 ) <= hist811 ( 31 downto 0 );
hist( 26015 downto 25984 ) <= hist812 ( 31 downto 0 );
hist( 26047 downto 26016 ) <= hist813 ( 31 downto 0 );
hist( 26079 downto 26048 ) <= hist814 ( 31 downto 0 );
hist( 26111 downto 26080 ) <= hist815 ( 31 downto 0 );
hist( 26143 downto 26112 ) <= hist816 ( 31 downto 0 );
hist( 26175 downto 26144 ) <= hist817 ( 31 downto 0 );
hist( 26207 downto 26176 ) <= hist818 ( 31 downto 0 );
hist( 26239 downto 26208 ) <= hist819 ( 31 downto 0 );
hist( 26271 downto 26240 ) <= hist820 ( 31 downto 0 );
hist( 26303 downto 26272 ) <= hist821 ( 31 downto 0 );
hist( 26335 downto 26304 ) <= hist822 ( 31 downto 0 );
hist( 26367 downto 26336 ) <= hist823 ( 31 downto 0 );
hist( 26399 downto 26368 ) <= hist824 ( 31 downto 0 );
hist( 26431 downto 26400 ) <= hist825 ( 31 downto 0 );
hist( 26463 downto 26432 ) <= hist826 ( 31 downto 0 );
hist( 26495 downto 26464 ) <= hist827 ( 31 downto 0 );
hist( 26527 downto 26496 ) <= hist828 ( 31 downto 0 );
hist( 26559 downto 26528 ) <= hist829 ( 31 downto 0 );
hist( 26591 downto 26560 ) <= hist830 ( 31 downto 0 );
hist( 26623 downto 26592 ) <= hist831 ( 31 downto 0 );
hist( 26655 downto 26624 ) <= hist832 ( 31 downto 0 );
hist( 26687 downto 26656 ) <= hist833 ( 31 downto 0 );
hist( 26719 downto 26688 ) <= hist834 ( 31 downto 0 );
hist( 26751 downto 26720 ) <= hist835 ( 31 downto 0 );
hist( 26783 downto 26752 ) <= hist836 ( 31 downto 0 );
hist( 26815 downto 26784 ) <= hist837 ( 31 downto 0 );
hist( 26847 downto 26816 ) <= hist838 ( 31 downto 0 );
hist( 26879 downto 26848 ) <= hist839 ( 31 downto 0 );
hist( 26911 downto 26880 ) <= hist840 ( 31 downto 0 );
hist( 26943 downto 26912 ) <= hist841 ( 31 downto 0 );
hist( 26975 downto 26944 ) <= hist842 ( 31 downto 0 );
hist( 27007 downto 26976 ) <= hist843 ( 31 downto 0 );
hist( 27039 downto 27008 ) <= hist844 ( 31 downto 0 );
hist( 27071 downto 27040 ) <= hist845 ( 31 downto 0 );
hist( 27103 downto 27072 ) <= hist846 ( 31 downto 0 );
hist( 27135 downto 27104 ) <= hist847 ( 31 downto 0 );
hist( 27167 downto 27136 ) <= hist848 ( 31 downto 0 );
hist( 27199 downto 27168 ) <= hist849 ( 31 downto 0 );
hist( 27231 downto 27200 ) <= hist850 ( 31 downto 0 );
hist( 27263 downto 27232 ) <= hist851 ( 31 downto 0 );
hist( 27295 downto 27264 ) <= hist852 ( 31 downto 0 );
hist( 27327 downto 27296 ) <= hist853 ( 31 downto 0 );
hist( 27359 downto 27328 ) <= hist854 ( 31 downto 0 );
hist( 27391 downto 27360 ) <= hist855 ( 31 downto 0 );
hist( 27423 downto 27392 ) <= hist856 ( 31 downto 0 );
hist( 27455 downto 27424 ) <= hist857 ( 31 downto 0 );
hist( 27487 downto 27456 ) <= hist858 ( 31 downto 0 );
hist( 27519 downto 27488 ) <= hist859 ( 31 downto 0 );
hist( 27551 downto 27520 ) <= hist860 ( 31 downto 0 );
hist( 27583 downto 27552 ) <= hist861 ( 31 downto 0 );
hist( 27615 downto 27584 ) <= hist862 ( 31 downto 0 );
hist( 27647 downto 27616 ) <= hist863 ( 31 downto 0 );
hist( 27679 downto 27648 ) <= hist864 ( 31 downto 0 );
hist( 27711 downto 27680 ) <= hist865 ( 31 downto 0 );
hist( 27743 downto 27712 ) <= hist866 ( 31 downto 0 );
hist( 27775 downto 27744 ) <= hist867 ( 31 downto 0 );
hist( 27807 downto 27776 ) <= hist868 ( 31 downto 0 );
hist( 27839 downto 27808 ) <= hist869 ( 31 downto 0 );
hist( 27871 downto 27840 ) <= hist870 ( 31 downto 0 );
hist( 27903 downto 27872 ) <= hist871 ( 31 downto 0 );
hist( 27935 downto 27904 ) <= hist872 ( 31 downto 0 );
hist( 27967 downto 27936 ) <= hist873 ( 31 downto 0 );
hist( 27999 downto 27968 ) <= hist874 ( 31 downto 0 );
hist( 28031 downto 28000 ) <= hist875 ( 31 downto 0 );
hist( 28063 downto 28032 ) <= hist876 ( 31 downto 0 );
hist( 28095 downto 28064 ) <= hist877 ( 31 downto 0 );
hist( 28127 downto 28096 ) <= hist878 ( 31 downto 0 );
hist( 28159 downto 28128 ) <= hist879 ( 31 downto 0 );
hist( 28191 downto 28160 ) <= hist880 ( 31 downto 0 );
hist( 28223 downto 28192 ) <= hist881 ( 31 downto 0 );
hist( 28255 downto 28224 ) <= hist882 ( 31 downto 0 );
hist( 28287 downto 28256 ) <= hist883 ( 31 downto 0 );
hist( 28319 downto 28288 ) <= hist884 ( 31 downto 0 );
hist( 28351 downto 28320 ) <= hist885 ( 31 downto 0 );
hist( 28383 downto 28352 ) <= hist886 ( 31 downto 0 );
hist( 28415 downto 28384 ) <= hist887 ( 31 downto 0 );
hist( 28447 downto 28416 ) <= hist888 ( 31 downto 0 );
hist( 28479 downto 28448 ) <= hist889 ( 31 downto 0 );
hist( 28511 downto 28480 ) <= hist890 ( 31 downto 0 );
hist( 28543 downto 28512 ) <= hist891 ( 31 downto 0 );
hist( 28575 downto 28544 ) <= hist892 ( 31 downto 0 );
hist( 28607 downto 28576 ) <= hist893 ( 31 downto 0 );
hist( 28639 downto 28608 ) <= hist894 ( 31 downto 0 );
hist( 28671 downto 28640 ) <= hist895 ( 31 downto 0 );
hist( 28703 downto 28672 ) <= hist896 ( 31 downto 0 );
hist( 28735 downto 28704 ) <= hist897 ( 31 downto 0 );
hist( 28767 downto 28736 ) <= hist898 ( 31 downto 0 );
hist( 28799 downto 28768 ) <= hist899 ( 31 downto 0 );
hist( 28831 downto 28800 ) <= hist900 ( 31 downto 0 );
hist( 28863 downto 28832 ) <= hist901 ( 31 downto 0 );
hist( 28895 downto 28864 ) <= hist902 ( 31 downto 0 );
hist( 28927 downto 28896 ) <= hist903 ( 31 downto 0 );
hist( 28959 downto 28928 ) <= hist904 ( 31 downto 0 );
hist( 28991 downto 28960 ) <= hist905 ( 31 downto 0 );
hist( 29023 downto 28992 ) <= hist906 ( 31 downto 0 );
hist( 29055 downto 29024 ) <= hist907 ( 31 downto 0 );
hist( 29087 downto 29056 ) <= hist908 ( 31 downto 0 );
hist( 29119 downto 29088 ) <= hist909 ( 31 downto 0 );
hist( 29151 downto 29120 ) <= hist910 ( 31 downto 0 );
hist( 29183 downto 29152 ) <= hist911 ( 31 downto 0 );
hist( 29215 downto 29184 ) <= hist912 ( 31 downto 0 );
hist( 29247 downto 29216 ) <= hist913 ( 31 downto 0 );
hist( 29279 downto 29248 ) <= hist914 ( 31 downto 0 );
hist( 29311 downto 29280 ) <= hist915 ( 31 downto 0 );
hist( 29343 downto 29312 ) <= hist916 ( 31 downto 0 );
hist( 29375 downto 29344 ) <= hist917 ( 31 downto 0 );
hist( 29407 downto 29376 ) <= hist918 ( 31 downto 0 );
hist( 29439 downto 29408 ) <= hist919 ( 31 downto 0 );
hist( 29471 downto 29440 ) <= hist920 ( 31 downto 0 );
hist( 29503 downto 29472 ) <= hist921 ( 31 downto 0 );
hist( 29535 downto 29504 ) <= hist922 ( 31 downto 0 );
hist( 29567 downto 29536 ) <= hist923 ( 31 downto 0 );
hist( 29599 downto 29568 ) <= hist924 ( 31 downto 0 );
hist( 29631 downto 29600 ) <= hist925 ( 31 downto 0 );
hist( 29663 downto 29632 ) <= hist926 ( 31 downto 0 );
hist( 29695 downto 29664 ) <= hist927 ( 31 downto 0 );
hist( 29727 downto 29696 ) <= hist928 ( 31 downto 0 );
hist( 29759 downto 29728 ) <= hist929 ( 31 downto 0 );
hist( 29791 downto 29760 ) <= hist930 ( 31 downto 0 );
hist( 29823 downto 29792 ) <= hist931 ( 31 downto 0 );
hist( 29855 downto 29824 ) <= hist932 ( 31 downto 0 );
hist( 29887 downto 29856 ) <= hist933 ( 31 downto 0 );
hist( 29919 downto 29888 ) <= hist934 ( 31 downto 0 );
hist( 29951 downto 29920 ) <= hist935 ( 31 downto 0 );
hist( 29983 downto 29952 ) <= hist936 ( 31 downto 0 );
hist( 30015 downto 29984 ) <= hist937 ( 31 downto 0 );
hist( 30047 downto 30016 ) <= hist938 ( 31 downto 0 );
hist( 30079 downto 30048 ) <= hist939 ( 31 downto 0 );
hist( 30111 downto 30080 ) <= hist940 ( 31 downto 0 );
hist( 30143 downto 30112 ) <= hist941 ( 31 downto 0 );
hist( 30175 downto 30144 ) <= hist942 ( 31 downto 0 );
hist( 30207 downto 30176 ) <= hist943 ( 31 downto 0 );
hist( 30239 downto 30208 ) <= hist944 ( 31 downto 0 );
hist( 30271 downto 30240 ) <= hist945 ( 31 downto 0 );
hist( 30303 downto 30272 ) <= hist946 ( 31 downto 0 );
hist( 30335 downto 30304 ) <= hist947 ( 31 downto 0 );
hist( 30367 downto 30336 ) <= hist948 ( 31 downto 0 );
hist( 30399 downto 30368 ) <= hist949 ( 31 downto 0 );
hist( 30431 downto 30400 ) <= hist950 ( 31 downto 0 );
hist( 30463 downto 30432 ) <= hist951 ( 31 downto 0 );
hist( 30495 downto 30464 ) <= hist952 ( 31 downto 0 );
hist( 30527 downto 30496 ) <= hist953 ( 31 downto 0 );
hist( 30559 downto 30528 ) <= hist954 ( 31 downto 0 );
hist( 30591 downto 30560 ) <= hist955 ( 31 downto 0 );
hist( 30623 downto 30592 ) <= hist956 ( 31 downto 0 );
hist( 30655 downto 30624 ) <= hist957 ( 31 downto 0 );
hist( 30687 downto 30656 ) <= hist958 ( 31 downto 0 );
hist( 30719 downto 30688 ) <= hist959 ( 31 downto 0 );
hist( 30751 downto 30720 ) <= hist960 ( 31 downto 0 );
hist( 30783 downto 30752 ) <= hist961 ( 31 downto 0 );
hist( 30815 downto 30784 ) <= hist962 ( 31 downto 0 );
hist( 30847 downto 30816 ) <= hist963 ( 31 downto 0 );
hist( 30879 downto 30848 ) <= hist964 ( 31 downto 0 );
hist( 30911 downto 30880 ) <= hist965 ( 31 downto 0 );
hist( 30943 downto 30912 ) <= hist966 ( 31 downto 0 );
hist( 30975 downto 30944 ) <= hist967 ( 31 downto 0 );
hist( 31007 downto 30976 ) <= hist968 ( 31 downto 0 );
hist( 31039 downto 31008 ) <= hist969 ( 31 downto 0 );
hist( 31071 downto 31040 ) <= hist970 ( 31 downto 0 );
hist( 31103 downto 31072 ) <= hist971 ( 31 downto 0 );
hist( 31135 downto 31104 ) <= hist972 ( 31 downto 0 );
hist( 31167 downto 31136 ) <= hist973 ( 31 downto 0 );
hist( 31199 downto 31168 ) <= hist974 ( 31 downto 0 );
hist( 31231 downto 31200 ) <= hist975 ( 31 downto 0 );
hist( 31263 downto 31232 ) <= hist976 ( 31 downto 0 );
hist( 31295 downto 31264 ) <= hist977 ( 31 downto 0 );
hist( 31327 downto 31296 ) <= hist978 ( 31 downto 0 );
hist( 31359 downto 31328 ) <= hist979 ( 31 downto 0 );
hist( 31391 downto 31360 ) <= hist980 ( 31 downto 0 );
hist( 31423 downto 31392 ) <= hist981 ( 31 downto 0 );
hist( 31455 downto 31424 ) <= hist982 ( 31 downto 0 );
hist( 31487 downto 31456 ) <= hist983 ( 31 downto 0 );
hist( 31519 downto 31488 ) <= hist984 ( 31 downto 0 );
hist( 31551 downto 31520 ) <= hist985 ( 31 downto 0 );
hist( 31583 downto 31552 ) <= hist986 ( 31 downto 0 );
hist( 31615 downto 31584 ) <= hist987 ( 31 downto 0 );
hist( 31647 downto 31616 ) <= hist988 ( 31 downto 0 );
hist( 31679 downto 31648 ) <= hist989 ( 31 downto 0 );
hist( 31711 downto 31680 ) <= hist990 ( 31 downto 0 );
hist( 31743 downto 31712 ) <= hist991 ( 31 downto 0 );
hist( 31775 downto 31744 ) <= hist992 ( 31 downto 0 );
hist( 31807 downto 31776 ) <= hist993 ( 31 downto 0 );
hist( 31839 downto 31808 ) <= hist994 ( 31 downto 0 );
hist( 31871 downto 31840 ) <= hist995 ( 31 downto 0 );
hist( 31903 downto 31872 ) <= hist996 ( 31 downto 0 );
hist( 31935 downto 31904 ) <= hist997 ( 31 downto 0 );
hist( 31967 downto 31936 ) <= hist998 ( 31 downto 0 );
hist( 31999 downto 31968 ) <= hist999 ( 31 downto 0 );
hist( 32031 downto 32000 ) <= hist1000 ( 31 downto 0 );
hist( 32063 downto 32032 ) <= hist1001 ( 31 downto 0 );
hist( 32095 downto 32064 ) <= hist1002 ( 31 downto 0 );
hist( 32127 downto 32096 ) <= hist1003 ( 31 downto 0 );
hist( 32159 downto 32128 ) <= hist1004 ( 31 downto 0 );
hist( 32191 downto 32160 ) <= hist1005 ( 31 downto 0 );
hist( 32223 downto 32192 ) <= hist1006 ( 31 downto 0 );
hist( 32255 downto 32224 ) <= hist1007 ( 31 downto 0 );
hist( 32287 downto 32256 ) <= hist1008 ( 31 downto 0 );
hist( 32319 downto 32288 ) <= hist1009 ( 31 downto 0 );
hist( 32351 downto 32320 ) <= hist1010 ( 31 downto 0 );
hist( 32383 downto 32352 ) <= hist1011 ( 31 downto 0 );
hist( 32415 downto 32384 ) <= hist1012 ( 31 downto 0 );
hist( 32447 downto 32416 ) <= hist1013 ( 31 downto 0 );
hist( 32479 downto 32448 ) <= hist1014 ( 31 downto 0 );
hist( 32511 downto 32480 ) <= hist1015 ( 31 downto 0 );
hist( 32543 downto 32512 ) <= hist1016 ( 31 downto 0 );
hist( 32575 downto 32544 ) <= hist1017 ( 31 downto 0 );
hist( 32607 downto 32576 ) <= hist1018 ( 31 downto 0 );
hist( 32639 downto 32608 ) <= hist1019 ( 31 downto 0 );
hist( 32671 downto 32640 ) <= hist1020 ( 31 downto 0 );
hist( 32703 downto 32672 ) <= hist1021 ( 31 downto 0 );
hist( 32735 downto 32704 ) <= hist1022 ( 31 downto 0 );
hist( 32767 downto 32736 ) <= hist1023 ( 31 downto 0 );

total_time <= time_gone;

Pout <= out_tmp;

end Behavioral;

